-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbb",
     9 => x"c0080b0b",
    10 => x"0bbbc408",
    11 => x"0b0b0bbb",
    12 => x"c8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bbc80c0b",
    16 => x"0b0bbbc4",
    17 => x"0c0b0b0b",
    18 => x"bbc00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb194",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bbc07080",
    57 => x"c5f0278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188c504",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbbd00c",
    65 => x"9f0bbbd4",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bbd408ff",
    69 => x"05bbd40c",
    70 => x"bbd40880",
    71 => x"25eb38bb",
    72 => x"d008ff05",
    73 => x"bbd00cbb",
    74 => x"d0088025",
    75 => x"d738800b",
    76 => x"bbd40c80",
    77 => x"0bbbd00c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbbd008",
    97 => x"258f3882",
    98 => x"bd2dbbd0",
    99 => x"08ff05bb",
   100 => x"d00c82ff",
   101 => x"04bbd008",
   102 => x"bbd40853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bbd008a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134bbd4",
   111 => x"088105bb",
   112 => x"d40cbbd4",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbbd40c",
   116 => x"bbd00881",
   117 => x"05bbd00c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134bb",
   122 => x"d4088105",
   123 => x"bbd40cbb",
   124 => x"d408a02e",
   125 => x"0981068e",
   126 => x"38800bbb",
   127 => x"d40cbbd0",
   128 => x"088105bb",
   129 => x"d00c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbbd8",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbbd80c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872bb",
   169 => x"d8088407",
   170 => x"bbd80c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb6fc",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"bbd80852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bbc00c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"92710c86",
   219 => x"a42d8271",
   220 => x"0c028405",
   221 => x"0d0402dc",
   222 => x"050d7a54",
   223 => x"807453bb",
   224 => x"dc5259a8",
   225 => x"b32dbbc0",
   226 => x"08792e81",
   227 => x"9138bbe0",
   228 => x"0870f80c",
   229 => x"891580f5",
   230 => x"2d8a1680",
   231 => x"f52d7182",
   232 => x"80290588",
   233 => x"1780f52d",
   234 => x"70848080",
   235 => x"2912f40c",
   236 => x"57555755",
   237 => x"a40bec0c",
   238 => x"78ff1655",
   239 => x"5873792e",
   240 => x"8b388118",
   241 => x"74812a55",
   242 => x"5873f738",
   243 => x"f7185881",
   244 => x"59807525",
   245 => x"80c83877",
   246 => x"52735184",
   247 => x"8b2dbca8",
   248 => x"52bbdc51",
   249 => x"aaf22dbb",
   250 => x"c008802e",
   251 => x"9a38bca8",
   252 => x"5783fc56",
   253 => x"76708405",
   254 => x"5808e80c",
   255 => x"fc165675",
   256 => x"8025f138",
   257 => x"888e04bb",
   258 => x"c0085984",
   259 => x"8055bbdc",
   260 => x"51aac42d",
   261 => x"fc801581",
   262 => x"15555587",
   263 => x"d10486b7",
   264 => x"2d840bec",
   265 => x"0c78802e",
   266 => x"8d38b780",
   267 => x"5190dd2d",
   268 => x"8ee02d88",
   269 => x"bc04b990",
   270 => x"5190dd2d",
   271 => x"78bbc00c",
   272 => x"02a4050d",
   273 => x"0402e005",
   274 => x"0d805584",
   275 => x"0bec0c8e",
   276 => x"c12d8bab",
   277 => x"2d81f82d",
   278 => x"9fac2dbb",
   279 => x"c008752e",
   280 => x"82b4388c",
   281 => x"0bec0cb5",
   282 => x"bc52bbdc",
   283 => x"51a8b32d",
   284 => x"bbc00875",
   285 => x"2e80e538",
   286 => x"bbe00875",
   287 => x"ff125659",
   288 => x"5673752e",
   289 => x"8b388118",
   290 => x"74812a55",
   291 => x"5873f738",
   292 => x"f7185880",
   293 => x"762580c4",
   294 => x"38775273",
   295 => x"51848b2d",
   296 => x"bca852bb",
   297 => x"dc51aaf2",
   298 => x"2dbbc008",
   299 => x"802e9a38",
   300 => x"bca85783",
   301 => x"fc557670",
   302 => x"84055808",
   303 => x"e80cfc15",
   304 => x"55748025",
   305 => x"f13889cc",
   306 => x"04848056",
   307 => x"bbdc51aa",
   308 => x"c42dfc80",
   309 => x"16811555",
   310 => x"56899304",
   311 => x"bbe008f8",
   312 => x"0c86b72d",
   313 => x"840bec0c",
   314 => x"86f651b1",
   315 => x"8c2db780",
   316 => x"5190dd2d",
   317 => x"8ee02d8b",
   318 => x"b72d90ed",
   319 => x"2db7a00b",
   320 => x"80f52d70",
   321 => x"822b8c06",
   322 => x"b7940b80",
   323 => x"f52d8306",
   324 => x"7107b7ac",
   325 => x"0b80f52d",
   326 => x"70842bb0",
   327 => x"06b7b80b",
   328 => x"80f52d70",
   329 => x"862b81c0",
   330 => x"06747307",
   331 => x"07b7c40b",
   332 => x"80f52d70",
   333 => x"882b8280",
   334 => x"06b7d00b",
   335 => x"80f52d70",
   336 => x"892b8480",
   337 => x"06747307",
   338 => x"07b7dc0b",
   339 => x"80f52d70",
   340 => x"8a2b9880",
   341 => x"06b7e80b",
   342 => x"80f52d70",
   343 => x"8c2b81e0",
   344 => x"80067473",
   345 => x"0707b7f4",
   346 => x"0b80f52d",
   347 => x"708f2b82",
   348 => x"80800672",
   349 => x"07fc0c53",
   350 => x"54545454",
   351 => x"54545454",
   352 => x"545b5452",
   353 => x"57545486",
   354 => x"53bbc008",
   355 => x"83388453",
   356 => x"72ec0c89",
   357 => x"f704800b",
   358 => x"bbc00c02",
   359 => x"a0050d04",
   360 => x"71980c04",
   361 => x"ffb008bb",
   362 => x"c00c0481",
   363 => x"0bffb00c",
   364 => x"04800bff",
   365 => x"b00c0402",
   366 => x"f4050d8c",
   367 => x"b904bbc0",
   368 => x"0881f02e",
   369 => x"09810689",
   370 => x"38810bb9",
   371 => x"f40c8cb9",
   372 => x"04bbc008",
   373 => x"81e02e09",
   374 => x"81068938",
   375 => x"810bb9f8",
   376 => x"0c8cb904",
   377 => x"bbc00852",
   378 => x"b9f80880",
   379 => x"2e8838bb",
   380 => x"c0088180",
   381 => x"05527184",
   382 => x"2c728f06",
   383 => x"5353b9f4",
   384 => x"08802e99",
   385 => x"38728429",
   386 => x"b9b40572",
   387 => x"1381712b",
   388 => x"70097308",
   389 => x"06730c51",
   390 => x"53538caf",
   391 => x"04728429",
   392 => x"b9b40572",
   393 => x"1383712b",
   394 => x"72080772",
   395 => x"0c535380",
   396 => x"0bb9f80c",
   397 => x"800bb9f4",
   398 => x"0cbbe851",
   399 => x"8dba2dbb",
   400 => x"c008ff24",
   401 => x"fef83880",
   402 => x"0bbbc00c",
   403 => x"028c050d",
   404 => x"0402f805",
   405 => x"0db9b452",
   406 => x"8f518072",
   407 => x"70840554",
   408 => x"0cff1151",
   409 => x"708025f2",
   410 => x"38028805",
   411 => x"0d0402f0",
   412 => x"050d7551",
   413 => x"8bb12d70",
   414 => x"822cfc06",
   415 => x"b9b41172",
   416 => x"109e0671",
   417 => x"0870722a",
   418 => x"70830682",
   419 => x"742b7009",
   420 => x"7406760c",
   421 => x"54515657",
   422 => x"5351538b",
   423 => x"ab2d71bb",
   424 => x"c00c0290",
   425 => x"050d0402",
   426 => x"fc050d72",
   427 => x"5180710c",
   428 => x"800b8412",
   429 => x"0c028405",
   430 => x"0d0402f0",
   431 => x"050d7570",
   432 => x"08841208",
   433 => x"535353ff",
   434 => x"5471712e",
   435 => x"a8388bb1",
   436 => x"2d841308",
   437 => x"70842914",
   438 => x"88117008",
   439 => x"7081ff06",
   440 => x"84180881",
   441 => x"11870684",
   442 => x"1a0c5351",
   443 => x"55515151",
   444 => x"8bab2d71",
   445 => x"5473bbc0",
   446 => x"0c029005",
   447 => x"0d0402f8",
   448 => x"050d8bb1",
   449 => x"2de00870",
   450 => x"8b2a7081",
   451 => x"06515252",
   452 => x"70802e9d",
   453 => x"38bbe808",
   454 => x"708429bb",
   455 => x"f0057381",
   456 => x"ff06710c",
   457 => x"5151bbe8",
   458 => x"08811187",
   459 => x"06bbe80c",
   460 => x"51800bbc",
   461 => x"900c8ba4",
   462 => x"2d8bab2d",
   463 => x"0288050d",
   464 => x"0402fc05",
   465 => x"0dbbe851",
   466 => x"8da72d8c",
   467 => x"d12d8dfe",
   468 => x"518ba02d",
   469 => x"0284050d",
   470 => x"04bc9408",
   471 => x"bbc00c04",
   472 => x"02fc050d",
   473 => x"8eea048b",
   474 => x"b72d80f6",
   475 => x"518cee2d",
   476 => x"bbc008f3",
   477 => x"3880da51",
   478 => x"8cee2dbb",
   479 => x"c008e838",
   480 => x"bbc008ba",
   481 => x"800cbbc0",
   482 => x"085184f0",
   483 => x"2d028405",
   484 => x"0d0402ec",
   485 => x"050d7654",
   486 => x"8052870b",
   487 => x"881580f5",
   488 => x"2d565374",
   489 => x"72248338",
   490 => x"a0537251",
   491 => x"82f92d81",
   492 => x"128b1580",
   493 => x"f52d5452",
   494 => x"727225de",
   495 => x"38029405",
   496 => x"0d0402f0",
   497 => x"050dbc94",
   498 => x"085481f8",
   499 => x"2d800bbc",
   500 => x"980c7308",
   501 => x"802e8180",
   502 => x"38820bbb",
   503 => x"d40cbc98",
   504 => x"088f06bb",
   505 => x"d00c7308",
   506 => x"5271832e",
   507 => x"96387183",
   508 => x"26893871",
   509 => x"812eaf38",
   510 => x"90c30471",
   511 => x"852e9f38",
   512 => x"90c30488",
   513 => x"1480f52d",
   514 => x"841508b5",
   515 => x"c8535452",
   516 => x"85fe2d71",
   517 => x"84291370",
   518 => x"08525290",
   519 => x"c7047351",
   520 => x"8f922d90",
   521 => x"c304b9fc",
   522 => x"08881508",
   523 => x"2c708106",
   524 => x"51527180",
   525 => x"2e8738b5",
   526 => x"cc5190c0",
   527 => x"04b5d051",
   528 => x"85fe2d84",
   529 => x"14085185",
   530 => x"fe2dbc98",
   531 => x"088105bc",
   532 => x"980c8c14",
   533 => x"548fd204",
   534 => x"0290050d",
   535 => x"0471bc94",
   536 => x"0c8fc22d",
   537 => x"bc9808ff",
   538 => x"05bc9c0c",
   539 => x"0402e805",
   540 => x"0dbc9408",
   541 => x"bca00857",
   542 => x"5587518c",
   543 => x"ee2dbbc0",
   544 => x"08812a70",
   545 => x"81065152",
   546 => x"71802ea0",
   547 => x"38919304",
   548 => x"8bb72d87",
   549 => x"518cee2d",
   550 => x"bbc008f4",
   551 => x"38ba8008",
   552 => x"813270ba",
   553 => x"800c7052",
   554 => x"5284f02d",
   555 => x"80fe518c",
   556 => x"ee2dbbc0",
   557 => x"08802ea6",
   558 => x"38ba8008",
   559 => x"802e9138",
   560 => x"800bba80",
   561 => x"0c805184",
   562 => x"f02d91d0",
   563 => x"048bb72d",
   564 => x"80fe518c",
   565 => x"ee2dbbc0",
   566 => x"08f33886",
   567 => x"e22dba80",
   568 => x"08903881",
   569 => x"fd518cee",
   570 => x"2d81fa51",
   571 => x"8cee2d97",
   572 => x"a30481f5",
   573 => x"518cee2d",
   574 => x"bbc00881",
   575 => x"2a708106",
   576 => x"51527180",
   577 => x"2eaf38bc",
   578 => x"9c085271",
   579 => x"802e8938",
   580 => x"ff12bc9c",
   581 => x"0c92b504",
   582 => x"bc980810",
   583 => x"bc980805",
   584 => x"70842916",
   585 => x"51528812",
   586 => x"08802e89",
   587 => x"38ff5188",
   588 => x"12085271",
   589 => x"2d81f251",
   590 => x"8cee2dbb",
   591 => x"c008812a",
   592 => x"70810651",
   593 => x"5271802e",
   594 => x"b138bc98",
   595 => x"08ff11bc",
   596 => x"9c085653",
   597 => x"53737225",
   598 => x"89388114",
   599 => x"bc9c0c92",
   600 => x"fa047210",
   601 => x"13708429",
   602 => x"16515288",
   603 => x"1208802e",
   604 => x"8938fe51",
   605 => x"88120852",
   606 => x"712d81fd",
   607 => x"518cee2d",
   608 => x"bbc00881",
   609 => x"2a708106",
   610 => x"51527180",
   611 => x"2ead38bc",
   612 => x"9c08802e",
   613 => x"8938800b",
   614 => x"bc9c0c93",
   615 => x"bb04bc98",
   616 => x"0810bc98",
   617 => x"08057084",
   618 => x"29165152",
   619 => x"88120880",
   620 => x"2e8938fd",
   621 => x"51881208",
   622 => x"52712d81",
   623 => x"fa518cee",
   624 => x"2dbbc008",
   625 => x"812a7081",
   626 => x"06515271",
   627 => x"802eae38",
   628 => x"bc9808ff",
   629 => x"115452bc",
   630 => x"9c087325",
   631 => x"883872bc",
   632 => x"9c0c93fd",
   633 => x"04711012",
   634 => x"70842916",
   635 => x"51528812",
   636 => x"08802e89",
   637 => x"38fc5188",
   638 => x"12085271",
   639 => x"2dbc9c08",
   640 => x"70535473",
   641 => x"802e8a38",
   642 => x"8c15ff15",
   643 => x"55559483",
   644 => x"04820bbb",
   645 => x"d40c718f",
   646 => x"06bbd00c",
   647 => x"81eb518c",
   648 => x"ee2dbbc0",
   649 => x"08812a70",
   650 => x"81065152",
   651 => x"71802ead",
   652 => x"38740885",
   653 => x"2e098106",
   654 => x"a4388815",
   655 => x"80f52dff",
   656 => x"05527188",
   657 => x"1681b72d",
   658 => x"71982b52",
   659 => x"71802588",
   660 => x"38800b88",
   661 => x"1681b72d",
   662 => x"74518f92",
   663 => x"2d81f451",
   664 => x"8cee2dbb",
   665 => x"c008812a",
   666 => x"70810651",
   667 => x"5271802e",
   668 => x"b3387408",
   669 => x"852e0981",
   670 => x"06aa3888",
   671 => x"1580f52d",
   672 => x"81055271",
   673 => x"881681b7",
   674 => x"2d7181ff",
   675 => x"068b1680",
   676 => x"f52d5452",
   677 => x"72722787",
   678 => x"38728816",
   679 => x"81b72d74",
   680 => x"518f922d",
   681 => x"80da518c",
   682 => x"ee2dbbc0",
   683 => x"08812a70",
   684 => x"81065152",
   685 => x"71802e81",
   686 => x"a638bc94",
   687 => x"08bc9c08",
   688 => x"55537380",
   689 => x"2e8a388c",
   690 => x"13ff1555",
   691 => x"5395c204",
   692 => x"72085271",
   693 => x"822ea638",
   694 => x"71822689",
   695 => x"3871812e",
   696 => x"a93896df",
   697 => x"0471832e",
   698 => x"b1387184",
   699 => x"2e098106",
   700 => x"80ed3888",
   701 => x"13085190",
   702 => x"dd2d96df",
   703 => x"04bc9c08",
   704 => x"51881308",
   705 => x"52712d96",
   706 => x"df04810b",
   707 => x"8814082b",
   708 => x"b9fc0832",
   709 => x"b9fc0c96",
   710 => x"b5048813",
   711 => x"80f52d81",
   712 => x"058b1480",
   713 => x"f52d5354",
   714 => x"71742483",
   715 => x"38805473",
   716 => x"881481b7",
   717 => x"2d8fc22d",
   718 => x"96df0475",
   719 => x"08802ea2",
   720 => x"38750851",
   721 => x"8cee2dbb",
   722 => x"c0088106",
   723 => x"5271802e",
   724 => x"8b38bc9c",
   725 => x"08518416",
   726 => x"0852712d",
   727 => x"88165675",
   728 => x"da388054",
   729 => x"800bbbd4",
   730 => x"0c738f06",
   731 => x"bbd00ca0",
   732 => x"5273bc9c",
   733 => x"082e0981",
   734 => x"069838bc",
   735 => x"9808ff05",
   736 => x"74327009",
   737 => x"81057072",
   738 => x"079f2a91",
   739 => x"71315151",
   740 => x"53537151",
   741 => x"82f92d81",
   742 => x"14548e74",
   743 => x"25c638ba",
   744 => x"80085271",
   745 => x"bbc00c02",
   746 => x"98050d04",
   747 => x"02f4050d",
   748 => x"d45281ff",
   749 => x"720c7108",
   750 => x"5381ff72",
   751 => x"0c72882b",
   752 => x"83fe8006",
   753 => x"72087081",
   754 => x"ff065152",
   755 => x"5381ff72",
   756 => x"0c727107",
   757 => x"882b7208",
   758 => x"7081ff06",
   759 => x"51525381",
   760 => x"ff720c72",
   761 => x"7107882b",
   762 => x"72087081",
   763 => x"ff067207",
   764 => x"bbc00c52",
   765 => x"53028c05",
   766 => x"0d0402f4",
   767 => x"050d7476",
   768 => x"7181ff06",
   769 => x"d40c5353",
   770 => x"bca40885",
   771 => x"3871892b",
   772 => x"5271982a",
   773 => x"d40c7190",
   774 => x"2a7081ff",
   775 => x"06d40c51",
   776 => x"71882a70",
   777 => x"81ff06d4",
   778 => x"0c517181",
   779 => x"ff06d40c",
   780 => x"72902a70",
   781 => x"81ff06d4",
   782 => x"0c51d408",
   783 => x"7081ff06",
   784 => x"515182b8",
   785 => x"bf527081",
   786 => x"ff2e0981",
   787 => x"06943881",
   788 => x"ff0bd40c",
   789 => x"d4087081",
   790 => x"ff06ff14",
   791 => x"54515171",
   792 => x"e53870bb",
   793 => x"c00c028c",
   794 => x"050d0402",
   795 => x"fc050d81",
   796 => x"c75181ff",
   797 => x"0bd40cff",
   798 => x"11517080",
   799 => x"25f43802",
   800 => x"84050d04",
   801 => x"02f4050d",
   802 => x"81ff0bd4",
   803 => x"0c935380",
   804 => x"5287fc80",
   805 => x"c15197fa",
   806 => x"2dbbc008",
   807 => x"8b3881ff",
   808 => x"0bd40c81",
   809 => x"5399b104",
   810 => x"98eb2dff",
   811 => x"135372df",
   812 => x"3872bbc0",
   813 => x"0c028c05",
   814 => x"0d0402ec",
   815 => x"050d810b",
   816 => x"bca40c84",
   817 => x"54d00870",
   818 => x"8f2a7081",
   819 => x"06515153",
   820 => x"72f33872",
   821 => x"d00c98eb",
   822 => x"2db5d451",
   823 => x"85fe2dd0",
   824 => x"08708f2a",
   825 => x"70810651",
   826 => x"515372f3",
   827 => x"38810bd0",
   828 => x"0cb15380",
   829 => x"5284d480",
   830 => x"c05197fa",
   831 => x"2dbbc008",
   832 => x"812e9338",
   833 => x"72822ebd",
   834 => x"38ff1353",
   835 => x"72e538ff",
   836 => x"145473ff",
   837 => x"b03898eb",
   838 => x"2d83aa52",
   839 => x"849c80c8",
   840 => x"5197fa2d",
   841 => x"bbc00881",
   842 => x"2e098106",
   843 => x"923897ac",
   844 => x"2dbbc008",
   845 => x"83ffff06",
   846 => x"537283aa",
   847 => x"2e9d3899",
   848 => x"842d9ad6",
   849 => x"04b5e051",
   850 => x"85fe2d80",
   851 => x"539ca404",
   852 => x"b5f85185",
   853 => x"fe2d8054",
   854 => x"9bf60481",
   855 => x"ff0bd40c",
   856 => x"b15498eb",
   857 => x"2d8fcf53",
   858 => x"805287fc",
   859 => x"80f75197",
   860 => x"fa2dbbc0",
   861 => x"0855bbc0",
   862 => x"08812e09",
   863 => x"81069b38",
   864 => x"81ff0bd4",
   865 => x"0c820a52",
   866 => x"849c80e9",
   867 => x"5197fa2d",
   868 => x"bbc00880",
   869 => x"2e8d3898",
   870 => x"eb2dff13",
   871 => x"5372c938",
   872 => x"9be90481",
   873 => x"ff0bd40c",
   874 => x"bbc00852",
   875 => x"87fc80fa",
   876 => x"5197fa2d",
   877 => x"bbc008b1",
   878 => x"3881ff0b",
   879 => x"d40cd408",
   880 => x"5381ff0b",
   881 => x"d40c81ff",
   882 => x"0bd40c81",
   883 => x"ff0bd40c",
   884 => x"81ff0bd4",
   885 => x"0c72862a",
   886 => x"70810676",
   887 => x"56515372",
   888 => x"9538bbc0",
   889 => x"08549bf6",
   890 => x"0473822e",
   891 => x"fee238ff",
   892 => x"145473fe",
   893 => x"ed3873bc",
   894 => x"a40c738b",
   895 => x"38815287",
   896 => x"fc80d051",
   897 => x"97fa2d81",
   898 => x"ff0bd40c",
   899 => x"d008708f",
   900 => x"2a708106",
   901 => x"51515372",
   902 => x"f33872d0",
   903 => x"0c81ff0b",
   904 => x"d40c8153",
   905 => x"72bbc00c",
   906 => x"0294050d",
   907 => x"0402e805",
   908 => x"0d785580",
   909 => x"5681ff0b",
   910 => x"d40cd008",
   911 => x"708f2a70",
   912 => x"81065151",
   913 => x"5372f338",
   914 => x"82810bd0",
   915 => x"0c81ff0b",
   916 => x"d40c7752",
   917 => x"87fc80d1",
   918 => x"5197fa2d",
   919 => x"80dbc6df",
   920 => x"54bbc008",
   921 => x"802e8a38",
   922 => x"b6985185",
   923 => x"fe2d9dc4",
   924 => x"0481ff0b",
   925 => x"d40cd408",
   926 => x"7081ff06",
   927 => x"51537281",
   928 => x"fe2e0981",
   929 => x"069d3880",
   930 => x"ff5397ac",
   931 => x"2dbbc008",
   932 => x"75708405",
   933 => x"570cff13",
   934 => x"53728025",
   935 => x"ed388156",
   936 => x"9da904ff",
   937 => x"145473c9",
   938 => x"3881ff0b",
   939 => x"d40c81ff",
   940 => x"0bd40cd0",
   941 => x"08708f2a",
   942 => x"70810651",
   943 => x"515372f3",
   944 => x"3872d00c",
   945 => x"75bbc00c",
   946 => x"0298050d",
   947 => x"0402e805",
   948 => x"0d77797b",
   949 => x"58555580",
   950 => x"53727625",
   951 => x"a3387470",
   952 => x"81055680",
   953 => x"f52d7470",
   954 => x"81055680",
   955 => x"f52d5252",
   956 => x"71712e86",
   957 => x"3881519e",
   958 => x"82048113",
   959 => x"539dd904",
   960 => x"805170bb",
   961 => x"c00c0298",
   962 => x"050d0402",
   963 => x"ec050d76",
   964 => x"5574802e",
   965 => x"be389a15",
   966 => x"80e02d51",
   967 => x"abcb2dbb",
   968 => x"c008bbc0",
   969 => x"0880c2d8",
   970 => x"0cbbc008",
   971 => x"545480c2",
   972 => x"b408802e",
   973 => x"99389415",
   974 => x"80e02d51",
   975 => x"abcb2dbb",
   976 => x"c008902b",
   977 => x"83fff00a",
   978 => x"06707507",
   979 => x"51537280",
   980 => x"c2d80c80",
   981 => x"c2d80853",
   982 => x"72802e9d",
   983 => x"3880c2ac",
   984 => x"08fe1471",
   985 => x"2980c2c0",
   986 => x"080580c2",
   987 => x"dc0c7084",
   988 => x"2b80c2b8",
   989 => x"0c549fa7",
   990 => x"0480c2c4",
   991 => x"0880c2d8",
   992 => x"0c80c2c8",
   993 => x"0880c2dc",
   994 => x"0c80c2b4",
   995 => x"08802e8b",
   996 => x"3880c2ac",
   997 => x"08842b53",
   998 => x"9fa20480",
   999 => x"c2cc0884",
  1000 => x"2b537280",
  1001 => x"c2b80c02",
  1002 => x"94050d04",
  1003 => x"02d8050d",
  1004 => x"800b80c2",
  1005 => x"b40c8454",
  1006 => x"99ba2dbb",
  1007 => x"c008802e",
  1008 => x"9538bca8",
  1009 => x"5280519c",
  1010 => x"ad2dbbc0",
  1011 => x"08802e86",
  1012 => x"38fe549f",
  1013 => x"de04ff14",
  1014 => x"54738024",
  1015 => x"db38738c",
  1016 => x"38b6a851",
  1017 => x"85fe2d73",
  1018 => x"55a58404",
  1019 => x"8056810b",
  1020 => x"80c2e00c",
  1021 => x"8853b6bc",
  1022 => x"52bcde51",
  1023 => x"9dcd2dbb",
  1024 => x"c008762e",
  1025 => x"09810688",
  1026 => x"38bbc008",
  1027 => x"80c2e00c",
  1028 => x"8853b6c8",
  1029 => x"52bcfa51",
  1030 => x"9dcd2dbb",
  1031 => x"c0088838",
  1032 => x"bbc00880",
  1033 => x"c2e00c80",
  1034 => x"c2e00880",
  1035 => x"2e80f838",
  1036 => x"bfee0b80",
  1037 => x"f52dbfef",
  1038 => x"0b80f52d",
  1039 => x"71982b71",
  1040 => x"902b07bf",
  1041 => x"f00b80f5",
  1042 => x"2d70882b",
  1043 => x"7207bff1",
  1044 => x"0b80f52d",
  1045 => x"710780c0",
  1046 => x"a60b80f5",
  1047 => x"2d80c0a7",
  1048 => x"0b80f52d",
  1049 => x"71882b07",
  1050 => x"535f5452",
  1051 => x"5a565755",
  1052 => x"7381abaa",
  1053 => x"2e098106",
  1054 => x"8d387551",
  1055 => x"ab9b2dbb",
  1056 => x"c00856a1",
  1057 => x"93047382",
  1058 => x"d4d52e87",
  1059 => x"38b6d451",
  1060 => x"a1d504bc",
  1061 => x"a8527551",
  1062 => x"9cad2dbb",
  1063 => x"c00855bb",
  1064 => x"c008802e",
  1065 => x"83de3888",
  1066 => x"53b6c852",
  1067 => x"bcfa519d",
  1068 => x"cd2dbbc0",
  1069 => x"088a3881",
  1070 => x"0b80c2b4",
  1071 => x"0ca1db04",
  1072 => x"8853b6bc",
  1073 => x"52bcde51",
  1074 => x"9dcd2dbb",
  1075 => x"c008802e",
  1076 => x"8a38b6e8",
  1077 => x"5185fe2d",
  1078 => x"a2b70480",
  1079 => x"c0a60b80",
  1080 => x"f52d5473",
  1081 => x"80d52e09",
  1082 => x"810680cb",
  1083 => x"3880c0a7",
  1084 => x"0b80f52d",
  1085 => x"547381aa",
  1086 => x"2e098106",
  1087 => x"ba38800b",
  1088 => x"bca80b80",
  1089 => x"f52d5654",
  1090 => x"7481e92e",
  1091 => x"83388154",
  1092 => x"7481eb2e",
  1093 => x"8c388055",
  1094 => x"73752e09",
  1095 => x"810682e4",
  1096 => x"38bcb30b",
  1097 => x"80f52d55",
  1098 => x"748d38bc",
  1099 => x"b40b80f5",
  1100 => x"2d547382",
  1101 => x"2e863880",
  1102 => x"55a58404",
  1103 => x"bcb50b80",
  1104 => x"f52d7080",
  1105 => x"c2ac0cff",
  1106 => x"0580c2b0",
  1107 => x"0cbcb60b",
  1108 => x"80f52dbc",
  1109 => x"b70b80f5",
  1110 => x"2d587605",
  1111 => x"77828029",
  1112 => x"057080c2",
  1113 => x"bc0cbcb8",
  1114 => x"0b80f52d",
  1115 => x"7080c2d0",
  1116 => x"0c80c2b4",
  1117 => x"08595758",
  1118 => x"76802e81",
  1119 => x"ac388853",
  1120 => x"b6c852bc",
  1121 => x"fa519dcd",
  1122 => x"2dbbc008",
  1123 => x"81f63880",
  1124 => x"c2ac0870",
  1125 => x"842b80c2",
  1126 => x"b80c7080",
  1127 => x"c2cc0cbc",
  1128 => x"cd0b80f5",
  1129 => x"2dbccc0b",
  1130 => x"80f52d71",
  1131 => x"82802905",
  1132 => x"bcce0b80",
  1133 => x"f52d7084",
  1134 => x"80802912",
  1135 => x"bccf0b80",
  1136 => x"f52d7081",
  1137 => x"800a2912",
  1138 => x"7080c2d4",
  1139 => x"0c80c2d0",
  1140 => x"08712980",
  1141 => x"c2bc0805",
  1142 => x"7080c2c0",
  1143 => x"0cbcd50b",
  1144 => x"80f52dbc",
  1145 => x"d40b80f5",
  1146 => x"2d718280",
  1147 => x"2905bcd6",
  1148 => x"0b80f52d",
  1149 => x"70848080",
  1150 => x"2912bcd7",
  1151 => x"0b80f52d",
  1152 => x"70982b81",
  1153 => x"f00a0672",
  1154 => x"057080c2",
  1155 => x"c40cfe11",
  1156 => x"7e297705",
  1157 => x"80c2c80c",
  1158 => x"52595243",
  1159 => x"545e5152",
  1160 => x"59525d57",
  1161 => x"5957a4fd",
  1162 => x"04bcba0b",
  1163 => x"80f52dbc",
  1164 => x"b90b80f5",
  1165 => x"2d718280",
  1166 => x"29057080",
  1167 => x"c2b80c70",
  1168 => x"a02983ff",
  1169 => x"0570892a",
  1170 => x"7080c2cc",
  1171 => x"0cbcbf0b",
  1172 => x"80f52dbc",
  1173 => x"be0b80f5",
  1174 => x"2d718280",
  1175 => x"29057080",
  1176 => x"c2d40c7b",
  1177 => x"71291e70",
  1178 => x"80c2c80c",
  1179 => x"7d80c2c4",
  1180 => x"0c730580",
  1181 => x"c2c00c55",
  1182 => x"5e515155",
  1183 => x"5580519e",
  1184 => x"8b2d8155",
  1185 => x"74bbc00c",
  1186 => x"02a8050d",
  1187 => x"0402ec05",
  1188 => x"0d767087",
  1189 => x"2c7180ff",
  1190 => x"06555654",
  1191 => x"80c2b408",
  1192 => x"8a387388",
  1193 => x"2c7481ff",
  1194 => x"065455bc",
  1195 => x"a85280c2",
  1196 => x"bc081551",
  1197 => x"9cad2dbb",
  1198 => x"c00854bb",
  1199 => x"c008802e",
  1200 => x"b43880c2",
  1201 => x"b408802e",
  1202 => x"98387284",
  1203 => x"29bca805",
  1204 => x"70085253",
  1205 => x"ab9b2dbb",
  1206 => x"c008f00a",
  1207 => x"0653a5f3",
  1208 => x"047210bc",
  1209 => x"a8057080",
  1210 => x"e02d5253",
  1211 => x"abcb2dbb",
  1212 => x"c0085372",
  1213 => x"5473bbc0",
  1214 => x"0c029405",
  1215 => x"0d0402e0",
  1216 => x"050d7970",
  1217 => x"842c80c2",
  1218 => x"dc080571",
  1219 => x"8f065255",
  1220 => x"53728938",
  1221 => x"bca85273",
  1222 => x"519cad2d",
  1223 => x"72a029bc",
  1224 => x"a8055480",
  1225 => x"7480f52d",
  1226 => x"56537473",
  1227 => x"2e833881",
  1228 => x"537481e5",
  1229 => x"2e81f138",
  1230 => x"81707406",
  1231 => x"54587280",
  1232 => x"2e81e538",
  1233 => x"8b1480f5",
  1234 => x"2d70832a",
  1235 => x"79065856",
  1236 => x"769938ba",
  1237 => x"84085372",
  1238 => x"89387280",
  1239 => x"c0a80b81",
  1240 => x"b72d76ba",
  1241 => x"840c7353",
  1242 => x"a8aa0475",
  1243 => x"8f2e0981",
  1244 => x"0681b538",
  1245 => x"749f068d",
  1246 => x"2980c09b",
  1247 => x"11515381",
  1248 => x"1480f52d",
  1249 => x"73708105",
  1250 => x"5581b72d",
  1251 => x"831480f5",
  1252 => x"2d737081",
  1253 => x"055581b7",
  1254 => x"2d851480",
  1255 => x"f52d7370",
  1256 => x"81055581",
  1257 => x"b72d8714",
  1258 => x"80f52d73",
  1259 => x"70810555",
  1260 => x"81b72d89",
  1261 => x"1480f52d",
  1262 => x"73708105",
  1263 => x"5581b72d",
  1264 => x"8e1480f5",
  1265 => x"2d737081",
  1266 => x"055581b7",
  1267 => x"2d901480",
  1268 => x"f52d7370",
  1269 => x"81055581",
  1270 => x"b72d9214",
  1271 => x"80f52d73",
  1272 => x"70810555",
  1273 => x"81b72d94",
  1274 => x"1480f52d",
  1275 => x"73708105",
  1276 => x"5581b72d",
  1277 => x"961480f5",
  1278 => x"2d737081",
  1279 => x"055581b7",
  1280 => x"2d981480",
  1281 => x"f52d7370",
  1282 => x"81055581",
  1283 => x"b72d9c14",
  1284 => x"80f52d73",
  1285 => x"70810555",
  1286 => x"81b72d9e",
  1287 => x"1480f52d",
  1288 => x"7381b72d",
  1289 => x"77ba840c",
  1290 => x"805372bb",
  1291 => x"c00c02a0",
  1292 => x"050d0402",
  1293 => x"cc050d7e",
  1294 => x"605e5a80",
  1295 => x"0b80c2d8",
  1296 => x"0880c2dc",
  1297 => x"08595c56",
  1298 => x"805880c2",
  1299 => x"b808782e",
  1300 => x"81b03877",
  1301 => x"8f06a017",
  1302 => x"5754738f",
  1303 => x"38bca852",
  1304 => x"76518117",
  1305 => x"579cad2d",
  1306 => x"bca85680",
  1307 => x"7680f52d",
  1308 => x"56547474",
  1309 => x"2e833881",
  1310 => x"547481e5",
  1311 => x"2e80f738",
  1312 => x"81707506",
  1313 => x"555c7380",
  1314 => x"2e80eb38",
  1315 => x"8b1680f5",
  1316 => x"2d980659",
  1317 => x"7880df38",
  1318 => x"8b537c52",
  1319 => x"75519dcd",
  1320 => x"2dbbc008",
  1321 => x"80d0389c",
  1322 => x"160851ab",
  1323 => x"9b2dbbc0",
  1324 => x"08841b0c",
  1325 => x"9a1680e0",
  1326 => x"2d51abcb",
  1327 => x"2dbbc008",
  1328 => x"bbc00888",
  1329 => x"1c0cbbc0",
  1330 => x"08555580",
  1331 => x"c2b40880",
  1332 => x"2e983894",
  1333 => x"1680e02d",
  1334 => x"51abcb2d",
  1335 => x"bbc00890",
  1336 => x"2b83fff0",
  1337 => x"0a067016",
  1338 => x"51547388",
  1339 => x"1b0c787a",
  1340 => x"0c7b54aa",
  1341 => x"bb048118",
  1342 => x"5880c2b8",
  1343 => x"087826fe",
  1344 => x"d23880c2",
  1345 => x"b408802e",
  1346 => x"b0387a51",
  1347 => x"a58d2dbb",
  1348 => x"c008bbc0",
  1349 => x"0880ffff",
  1350 => x"fff80655",
  1351 => x"5b7380ff",
  1352 => x"fffff82e",
  1353 => x"9438bbc0",
  1354 => x"08fe0580",
  1355 => x"c2ac0829",
  1356 => x"80c2c008",
  1357 => x"0557a8c8",
  1358 => x"04805473",
  1359 => x"bbc00c02",
  1360 => x"b4050d04",
  1361 => x"02f4050d",
  1362 => x"74700881",
  1363 => x"05710c70",
  1364 => x"0880c2b0",
  1365 => x"08065353",
  1366 => x"718e3888",
  1367 => x"130851a5",
  1368 => x"8d2dbbc0",
  1369 => x"0888140c",
  1370 => x"810bbbc0",
  1371 => x"0c028c05",
  1372 => x"0d0402f0",
  1373 => x"050d7588",
  1374 => x"1108fe05",
  1375 => x"80c2ac08",
  1376 => x"2980c2c0",
  1377 => x"08117208",
  1378 => x"80c2b008",
  1379 => x"06057955",
  1380 => x"5354549c",
  1381 => x"ad2d0290",
  1382 => x"050d0402",
  1383 => x"f4050d74",
  1384 => x"70882a83",
  1385 => x"fe800670",
  1386 => x"72982a07",
  1387 => x"72882b87",
  1388 => x"fc808006",
  1389 => x"73982b81",
  1390 => x"f00a0671",
  1391 => x"730707bb",
  1392 => x"c00c5651",
  1393 => x"5351028c",
  1394 => x"050d0402",
  1395 => x"f8050d02",
  1396 => x"8e0580f5",
  1397 => x"2d74882b",
  1398 => x"077083ff",
  1399 => x"ff06bbc0",
  1400 => x"0c510288",
  1401 => x"050d0402",
  1402 => x"f4050d74",
  1403 => x"76785354",
  1404 => x"52807125",
  1405 => x"97387270",
  1406 => x"81055480",
  1407 => x"f52d7270",
  1408 => x"81055481",
  1409 => x"b72dff11",
  1410 => x"5170eb38",
  1411 => x"807281b7",
  1412 => x"2d028c05",
  1413 => x"0d0402e8",
  1414 => x"050d7756",
  1415 => x"80705654",
  1416 => x"737624b3",
  1417 => x"3880c2b8",
  1418 => x"08742eab",
  1419 => x"387351a5",
  1420 => x"fe2dbbc0",
  1421 => x"08bbc008",
  1422 => x"09810570",
  1423 => x"bbc00807",
  1424 => x"9f2a7705",
  1425 => x"81175757",
  1426 => x"53537476",
  1427 => x"24893880",
  1428 => x"c2b80874",
  1429 => x"26d73872",
  1430 => x"bbc00c02",
  1431 => x"98050d04",
  1432 => x"02f0050d",
  1433 => x"bbbc0816",
  1434 => x"51ac962d",
  1435 => x"bbc00880",
  1436 => x"2e9e388b",
  1437 => x"53bbc008",
  1438 => x"5280c0a8",
  1439 => x"51abe72d",
  1440 => x"80c2e408",
  1441 => x"5473802e",
  1442 => x"873880c0",
  1443 => x"a851732d",
  1444 => x"0290050d",
  1445 => x"0402dc05",
  1446 => x"0d80705a",
  1447 => x"5574bbbc",
  1448 => x"0825b138",
  1449 => x"80c2b808",
  1450 => x"752ea938",
  1451 => x"7851a5fe",
  1452 => x"2dbbc008",
  1453 => x"09810570",
  1454 => x"bbc00807",
  1455 => x"9f2a7605",
  1456 => x"811b5b56",
  1457 => x"5474bbbc",
  1458 => x"08258938",
  1459 => x"80c2b808",
  1460 => x"7926d938",
  1461 => x"80557880",
  1462 => x"c2b80827",
  1463 => x"81d43878",
  1464 => x"51a5fe2d",
  1465 => x"bbc00880",
  1466 => x"2e81a838",
  1467 => x"bbc0088b",
  1468 => x"0580f52d",
  1469 => x"70842a70",
  1470 => x"81067710",
  1471 => x"78842b80",
  1472 => x"c0a80b80",
  1473 => x"f52d5c5c",
  1474 => x"53515556",
  1475 => x"73802e80",
  1476 => x"c9387416",
  1477 => x"822bafd6",
  1478 => x"0bba9012",
  1479 => x"0c547775",
  1480 => x"311080c2",
  1481 => x"e8115556",
  1482 => x"90747081",
  1483 => x"055681b7",
  1484 => x"2da07481",
  1485 => x"b72d7681",
  1486 => x"ff068116",
  1487 => x"58547380",
  1488 => x"2e8a389c",
  1489 => x"5380c0a8",
  1490 => x"52aed204",
  1491 => x"8b53bbc0",
  1492 => x"085280c2",
  1493 => x"ea1651af",
  1494 => x"8b047416",
  1495 => x"822bace0",
  1496 => x"0bba9012",
  1497 => x"0c547681",
  1498 => x"ff068116",
  1499 => x"58547380",
  1500 => x"2e8a389c",
  1501 => x"5380c0a8",
  1502 => x"52af8204",
  1503 => x"8b53bbc0",
  1504 => x"08527775",
  1505 => x"311080c2",
  1506 => x"e8055176",
  1507 => x"55abe72d",
  1508 => x"afa70474",
  1509 => x"90297531",
  1510 => x"701080c2",
  1511 => x"e8055154",
  1512 => x"bbc00874",
  1513 => x"81b72d81",
  1514 => x"1959748b",
  1515 => x"24a338ad",
  1516 => x"d6047490",
  1517 => x"29753170",
  1518 => x"1080c2e8",
  1519 => x"058c7731",
  1520 => x"57515480",
  1521 => x"7481b72d",
  1522 => x"9e14ff16",
  1523 => x"565474f3",
  1524 => x"3802a405",
  1525 => x"0d0402fc",
  1526 => x"050dbbbc",
  1527 => x"081351ac",
  1528 => x"962dbbc0",
  1529 => x"08802e88",
  1530 => x"38bbc008",
  1531 => x"519e8b2d",
  1532 => x"800bbbbc",
  1533 => x"0cad952d",
  1534 => x"8fc22d02",
  1535 => x"84050d04",
  1536 => x"02fc050d",
  1537 => x"725170fd",
  1538 => x"2ead3870",
  1539 => x"fd248a38",
  1540 => x"70fc2e80",
  1541 => x"c438b0e1",
  1542 => x"0470fe2e",
  1543 => x"b13870ff",
  1544 => x"2e098106",
  1545 => x"bc38bbbc",
  1546 => x"08517080",
  1547 => x"2eb338ff",
  1548 => x"11bbbc0c",
  1549 => x"b0e104bb",
  1550 => x"bc08f005",
  1551 => x"70bbbc0c",
  1552 => x"51708025",
  1553 => x"9c38800b",
  1554 => x"bbbc0cb0",
  1555 => x"e104bbbc",
  1556 => x"088105bb",
  1557 => x"bc0cb0e1",
  1558 => x"04bbbc08",
  1559 => x"9005bbbc",
  1560 => x"0cad952d",
  1561 => x"8fc22d02",
  1562 => x"84050d04",
  1563 => x"02fc050d",
  1564 => x"800bbbbc",
  1565 => x"0cad952d",
  1566 => x"8ed92dbb",
  1567 => x"c008bbac",
  1568 => x"0cba8851",
  1569 => x"90dd2d02",
  1570 => x"84050d04",
  1571 => x"7180c2e4",
  1572 => x"0c040000",
  1573 => x"00ffffff",
  1574 => x"ff00ffff",
  1575 => x"ffff00ff",
  1576 => x"ffffff00",
  1577 => x"52657365",
  1578 => x"74000000",
  1579 => x"43617267",
  1580 => x"61722044",
  1581 => x"6973636f",
  1582 => x"2f43696e",
  1583 => x"74612010",
  1584 => x"00000000",
  1585 => x"45786974",
  1586 => x"00000000",
  1587 => x"43617267",
  1588 => x"61206465",
  1589 => x"2043696e",
  1590 => x"74612052",
  1591 => x"61706964",
  1592 => x"61000000",
  1593 => x"43617267",
  1594 => x"61206465",
  1595 => x"2043696e",
  1596 => x"7461204e",
  1597 => x"6f726d61",
  1598 => x"6c000000",
  1599 => x"53706563",
  1600 => x"7472756d",
  1601 => x"20313238",
  1602 => x"4b000000",
  1603 => x"50656e74",
  1604 => x"61676f6e",
  1605 => x"20313032",
  1606 => x"344b0000",
  1607 => x"50726f66",
  1608 => x"69203130",
  1609 => x"32344b00",
  1610 => x"53706563",
  1611 => x"7472756d",
  1612 => x"2034384b",
  1613 => x"00000000",
  1614 => x"53706563",
  1615 => x"7472756d",
  1616 => x"202b3241",
  1617 => x"2f2b3300",
  1618 => x"554c412d",
  1619 => x"34380000",
  1620 => x"554c412d",
  1621 => x"31323800",
  1622 => x"50656e74",
  1623 => x"61676f6e",
  1624 => x"00000000",
  1625 => x"556c612b",
  1626 => x"20262054",
  1627 => x"696d6578",
  1628 => x"00000000",
  1629 => x"4e6f726d",
  1630 => x"616c0000",
  1631 => x"47656e65",
  1632 => x"72616c20",
  1633 => x"536f756e",
  1634 => x"6420324d",
  1635 => x"42000000",
  1636 => x"47656e65",
  1637 => x"72616c20",
  1638 => x"536f756e",
  1639 => x"64204465",
  1640 => x"73616374",
  1641 => x"69766164",
  1642 => x"6f000000",
  1643 => x"4d4d4320",
  1644 => x"43617264",
  1645 => x"206f6666",
  1646 => x"00000000",
  1647 => x"6469764d",
  1648 => x"4d430000",
  1649 => x"5a584d4d",
  1650 => x"43000000",
  1651 => x"4a6f7920",
  1652 => x"323a2053",
  1653 => x"696e636c",
  1654 => x"61697220",
  1655 => x"49000000",
  1656 => x"4a6f7920",
  1657 => x"323a2053",
  1658 => x"696e636c",
  1659 => x"61697220",
  1660 => x"49490000",
  1661 => x"4a6f7920",
  1662 => x"323a204b",
  1663 => x"656d7374",
  1664 => x"6f6e0000",
  1665 => x"4a6f7920",
  1666 => x"323a2043",
  1667 => x"7572736f",
  1668 => x"72000000",
  1669 => x"4a6f7920",
  1670 => x"313a2053",
  1671 => x"696e636c",
  1672 => x"61697220",
  1673 => x"49000000",
  1674 => x"4a6f7920",
  1675 => x"313a2053",
  1676 => x"696e636c",
  1677 => x"61697220",
  1678 => x"49490000",
  1679 => x"4a6f7920",
  1680 => x"313a204b",
  1681 => x"656d7374",
  1682 => x"6f6e0000",
  1683 => x"4a6f7920",
  1684 => x"313a2043",
  1685 => x"7572736f",
  1686 => x"72000000",
  1687 => x"5363616e",
  1688 => x"6c696e65",
  1689 => x"73204e6f",
  1690 => x"6e650000",
  1691 => x"5363616e",
  1692 => x"6c696e65",
  1693 => x"73204352",
  1694 => x"54203235",
  1695 => x"25000000",
  1696 => x"5363616e",
  1697 => x"6c696e65",
  1698 => x"73204352",
  1699 => x"54203530",
  1700 => x"25000000",
  1701 => x"5363616e",
  1702 => x"6c696e65",
  1703 => x"73204352",
  1704 => x"54203735",
  1705 => x"25000000",
  1706 => x"43617267",
  1707 => x"61204661",
  1708 => x"6c6c6964",
  1709 => x"61000000",
  1710 => x"4f4b0000",
  1711 => x"53504543",
  1712 => x"5452554d",
  1713 => x"44415400",
  1714 => x"16200000",
  1715 => x"14200000",
  1716 => x"15200000",
  1717 => x"53442069",
  1718 => x"6e69742e",
  1719 => x"2e2e0a00",
  1720 => x"53442063",
  1721 => x"61726420",
  1722 => x"72657365",
  1723 => x"74206661",
  1724 => x"696c6564",
  1725 => x"210a0000",
  1726 => x"53444843",
  1727 => x"20657272",
  1728 => x"6f72210a",
  1729 => x"00000000",
  1730 => x"57726974",
  1731 => x"65206661",
  1732 => x"696c6564",
  1733 => x"0a000000",
  1734 => x"52656164",
  1735 => x"20666169",
  1736 => x"6c65640a",
  1737 => x"00000000",
  1738 => x"43617264",
  1739 => x"20696e69",
  1740 => x"74206661",
  1741 => x"696c6564",
  1742 => x"0a000000",
  1743 => x"46415431",
  1744 => x"36202020",
  1745 => x"00000000",
  1746 => x"46415433",
  1747 => x"32202020",
  1748 => x"00000000",
  1749 => x"4e6f2070",
  1750 => x"61727469",
  1751 => x"74696f6e",
  1752 => x"20736967",
  1753 => x"0a000000",
  1754 => x"42616420",
  1755 => x"70617274",
  1756 => x"0a000000",
  1757 => x"4261636b",
  1758 => x"00000000",
  1759 => x"00000002",
  1760 => x"00000002",
  1761 => x"000018a4",
  1762 => x"0000034e",
  1763 => x"00000003",
  1764 => x"00001c80",
  1765 => x"00000004",
  1766 => x"00000003",
  1767 => x"00001c70",
  1768 => x"00000005",
  1769 => x"00000003",
  1770 => x"00001c60",
  1771 => x"00000005",
  1772 => x"00000003",
  1773 => x"00001c54",
  1774 => x"00000003",
  1775 => x"00000003",
  1776 => x"00001c4c",
  1777 => x"00000002",
  1778 => x"00000003",
  1779 => x"00001c44",
  1780 => x"00000002",
  1781 => x"00000003",
  1782 => x"00001c38",
  1783 => x"00000003",
  1784 => x"00000003",
  1785 => x"00001c24",
  1786 => x"00000005",
  1787 => x"00000003",
  1788 => x"00001c1c",
  1789 => x"00000002",
  1790 => x"00000002",
  1791 => x"000018ac",
  1792 => x"0000186c",
  1793 => x"00000002",
  1794 => x"000018c4",
  1795 => x"00000760",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"000018cc",
  1800 => x"000018e4",
  1801 => x"000018fc",
  1802 => x"0000190c",
  1803 => x"0000191c",
  1804 => x"00001928",
  1805 => x"00001938",
  1806 => x"00001948",
  1807 => x"00001950",
  1808 => x"00001958",
  1809 => x"00001964",
  1810 => x"00001974",
  1811 => x"0000197c",
  1812 => x"00001990",
  1813 => x"000019ac",
  1814 => x"000019bc",
  1815 => x"000019c4",
  1816 => x"000019cc",
  1817 => x"000019e0",
  1818 => x"000019f4",
  1819 => x"00001a04",
  1820 => x"00001a14",
  1821 => x"00001a28",
  1822 => x"00001a3c",
  1823 => x"00001a4c",
  1824 => x"00001a5c",
  1825 => x"00001a6c",
  1826 => x"00001a80",
  1827 => x"00001a94",
  1828 => x"00000004",
  1829 => x"00001aa8",
  1830 => x"00001c90",
  1831 => x"00000004",
  1832 => x"00001ab8",
  1833 => x"00001b80",
  1834 => x"00000000",
  1835 => x"00000000",
  1836 => x"00000000",
  1837 => x"00000000",
  1838 => x"00000000",
  1839 => x"00000000",
  1840 => x"00000000",
  1841 => x"00000000",
  1842 => x"00000000",
  1843 => x"00000000",
  1844 => x"00000000",
  1845 => x"00000000",
  1846 => x"00000000",
  1847 => x"00000000",
  1848 => x"00000000",
  1849 => x"00000000",
  1850 => x"00000000",
  1851 => x"00000000",
  1852 => x"00000000",
  1853 => x"00000000",
  1854 => x"00000000",
  1855 => x"00000000",
  1856 => x"00000000",
  1857 => x"00000000",
  1858 => x"00000002",
  1859 => x"00002168",
  1860 => x"00001660",
  1861 => x"00000002",
  1862 => x"00002186",
  1863 => x"00001660",
  1864 => x"00000002",
  1865 => x"000021a4",
  1866 => x"00001660",
  1867 => x"00000002",
  1868 => x"000021c2",
  1869 => x"00001660",
  1870 => x"00000002",
  1871 => x"000021e0",
  1872 => x"00001660",
  1873 => x"00000002",
  1874 => x"000021fe",
  1875 => x"00001660",
  1876 => x"00000002",
  1877 => x"0000221c",
  1878 => x"00001660",
  1879 => x"00000002",
  1880 => x"0000223a",
  1881 => x"00001660",
  1882 => x"00000002",
  1883 => x"00002258",
  1884 => x"00001660",
  1885 => x"00000002",
  1886 => x"00002276",
  1887 => x"00001660",
  1888 => x"00000002",
  1889 => x"00002294",
  1890 => x"00001660",
  1891 => x"00000002",
  1892 => x"000022b2",
  1893 => x"00001660",
  1894 => x"00000002",
  1895 => x"000022d0",
  1896 => x"00001660",
  1897 => x"00000004",
  1898 => x"00001b74",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00001800",
  1903 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

