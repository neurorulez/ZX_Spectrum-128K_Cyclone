-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbb",
     9 => x"c4080b0b",
    10 => x"0bbbc808",
    11 => x"0b0b0bbb",
    12 => x"cc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bbcc0c0b",
    16 => x"0b0bbbc8",
    17 => x"0c0b0b0b",
    18 => x"bbc40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb198",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bbc47080",
    57 => x"c5f4278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188c804",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbbd40c",
    65 => x"9f0bbbd8",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bbd808ff",
    69 => x"05bbd80c",
    70 => x"bbd80880",
    71 => x"25eb38bb",
    72 => x"d408ff05",
    73 => x"bbd40cbb",
    74 => x"d4088025",
    75 => x"d738800b",
    76 => x"bbd80c80",
    77 => x"0bbbd40c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbbd408",
    97 => x"258f3882",
    98 => x"bd2dbbd4",
    99 => x"08ff05bb",
   100 => x"d40c82ff",
   101 => x"04bbd408",
   102 => x"bbd80853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bbd408a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134bbd8",
   111 => x"088105bb",
   112 => x"d80cbbd8",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbbd80c",
   116 => x"bbd40881",
   117 => x"05bbd40c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134bb",
   122 => x"d8088105",
   123 => x"bbd80cbb",
   124 => x"d808a02e",
   125 => x"0981068e",
   126 => x"38800bbb",
   127 => x"d80cbbd4",
   128 => x"088105bb",
   129 => x"d40c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbbdc",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbbdc0c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872bb",
   169 => x"dc088407",
   170 => x"bbdc0c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb780",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"bbdc0852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bbc40c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"92710c86",
   219 => x"a42d8271",
   220 => x"0c028405",
   221 => x"0d0402dc",
   222 => x"050d7a54",
   223 => x"800bbbe4",
   224 => x"08f80c89",
   225 => x"1580f52d",
   226 => x"8a1680f5",
   227 => x"2d718280",
   228 => x"29058817",
   229 => x"80f52d70",
   230 => x"84808029",
   231 => x"12f40c52",
   232 => x"555659a4",
   233 => x"0bec0c73",
   234 => x"52bbe051",
   235 => x"a8b62dbb",
   236 => x"c408792e",
   237 => x"80eb38bb",
   238 => x"e40879ff",
   239 => x"12565956",
   240 => x"73792e8b",
   241 => x"38811874",
   242 => x"812a5558",
   243 => x"73f738f7",
   244 => x"18588159",
   245 => x"80762580",
   246 => x"c8387752",
   247 => x"7351848b",
   248 => x"2dbcac52",
   249 => x"bbe051aa",
   250 => x"f52dbbc4",
   251 => x"08802e9a",
   252 => x"38bcac57",
   253 => x"83fc5576",
   254 => x"70840558",
   255 => x"08e80cfc",
   256 => x"15557480",
   257 => x"25f13888",
   258 => x"9104bbc4",
   259 => x"08598480",
   260 => x"56bbe051",
   261 => x"aac72dfc",
   262 => x"80168115",
   263 => x"555687d4",
   264 => x"0486b72d",
   265 => x"840bec0c",
   266 => x"78802e8d",
   267 => x"38b78451",
   268 => x"90e02d8e",
   269 => x"e32d88bf",
   270 => x"04b99451",
   271 => x"90e02d78",
   272 => x"bbc40c02",
   273 => x"a4050d04",
   274 => x"02e0050d",
   275 => x"8055840b",
   276 => x"ec0c8ec4",
   277 => x"2d8bae2d",
   278 => x"81f82d9f",
   279 => x"af2dbbc4",
   280 => x"08752e82",
   281 => x"b4388c0b",
   282 => x"ec0cb5c0",
   283 => x"52bbe051",
   284 => x"a8b62dbb",
   285 => x"c408752e",
   286 => x"80e538bb",
   287 => x"e40875ff",
   288 => x"12565956",
   289 => x"73752e8b",
   290 => x"38811874",
   291 => x"812a5558",
   292 => x"73f738f7",
   293 => x"18588076",
   294 => x"2580c438",
   295 => x"77527351",
   296 => x"848b2dbc",
   297 => x"ac52bbe0",
   298 => x"51aaf52d",
   299 => x"bbc40880",
   300 => x"2e9a38bc",
   301 => x"ac5783fc",
   302 => x"55767084",
   303 => x"055808e8",
   304 => x"0cfc1555",
   305 => x"748025f1",
   306 => x"3889cf04",
   307 => x"848056bb",
   308 => x"e051aac7",
   309 => x"2dfc8016",
   310 => x"81155556",
   311 => x"899604bb",
   312 => x"e408f80c",
   313 => x"86b72d84",
   314 => x"0bec0c86",
   315 => x"f651b18f",
   316 => x"2db78451",
   317 => x"90e02d8e",
   318 => x"e32d8bba",
   319 => x"2d90f02d",
   320 => x"b7a40b80",
   321 => x"f52d7082",
   322 => x"2b8c06b7",
   323 => x"980b80f5",
   324 => x"2d830671",
   325 => x"07b7b00b",
   326 => x"80f52d70",
   327 => x"842bb006",
   328 => x"b7bc0b80",
   329 => x"f52d7086",
   330 => x"2b81c006",
   331 => x"74730707",
   332 => x"b7c80b80",
   333 => x"f52d7088",
   334 => x"2b828006",
   335 => x"b7d40b80",
   336 => x"f52d7089",
   337 => x"2b848006",
   338 => x"74730707",
   339 => x"b7e00b80",
   340 => x"f52d708a",
   341 => x"2b988006",
   342 => x"b7ec0b80",
   343 => x"f52d708c",
   344 => x"2b81e080",
   345 => x"06747307",
   346 => x"07b7f80b",
   347 => x"80f52d70",
   348 => x"8f2b8280",
   349 => x"80067207",
   350 => x"fc0c5354",
   351 => x"54545454",
   352 => x"54545454",
   353 => x"5b545257",
   354 => x"54548653",
   355 => x"bbc40883",
   356 => x"38845372",
   357 => x"ec0c89fa",
   358 => x"04800bbb",
   359 => x"c40c02a0",
   360 => x"050d0471",
   361 => x"980c04ff",
   362 => x"b008bbc4",
   363 => x"0c04810b",
   364 => x"ffb00c04",
   365 => x"800bffb0",
   366 => x"0c0402f4",
   367 => x"050d8cbc",
   368 => x"04bbc408",
   369 => x"81f02e09",
   370 => x"81068938",
   371 => x"810bb9f8",
   372 => x"0c8cbc04",
   373 => x"bbc40881",
   374 => x"e02e0981",
   375 => x"06893881",
   376 => x"0bb9fc0c",
   377 => x"8cbc04bb",
   378 => x"c40852b9",
   379 => x"fc08802e",
   380 => x"8838bbc4",
   381 => x"08818005",
   382 => x"5271842c",
   383 => x"728f0653",
   384 => x"53b9f808",
   385 => x"802e9938",
   386 => x"728429b9",
   387 => x"b8057213",
   388 => x"81712b70",
   389 => x"09730806",
   390 => x"730c5153",
   391 => x"538cb204",
   392 => x"728429b9",
   393 => x"b8057213",
   394 => x"83712b72",
   395 => x"0807720c",
   396 => x"5353800b",
   397 => x"b9fc0c80",
   398 => x"0bb9f80c",
   399 => x"bbec518d",
   400 => x"bd2dbbc4",
   401 => x"08ff24fe",
   402 => x"f838800b",
   403 => x"bbc40c02",
   404 => x"8c050d04",
   405 => x"02f8050d",
   406 => x"b9b8528f",
   407 => x"51807270",
   408 => x"8405540c",
   409 => x"ff115170",
   410 => x"8025f238",
   411 => x"0288050d",
   412 => x"0402f005",
   413 => x"0d75518b",
   414 => x"b42d7082",
   415 => x"2cfc06b9",
   416 => x"b8117210",
   417 => x"9e067108",
   418 => x"70722a70",
   419 => x"83068274",
   420 => x"2b700974",
   421 => x"06760c54",
   422 => x"51565753",
   423 => x"51538bae",
   424 => x"2d71bbc4",
   425 => x"0c029005",
   426 => x"0d0402fc",
   427 => x"050d7251",
   428 => x"80710c80",
   429 => x"0b84120c",
   430 => x"0284050d",
   431 => x"0402f005",
   432 => x"0d757008",
   433 => x"84120853",
   434 => x"5353ff54",
   435 => x"71712ea8",
   436 => x"388bb42d",
   437 => x"84130870",
   438 => x"84291488",
   439 => x"11700870",
   440 => x"81ff0684",
   441 => x"18088111",
   442 => x"8706841a",
   443 => x"0c535155",
   444 => x"5151518b",
   445 => x"ae2d7154",
   446 => x"73bbc40c",
   447 => x"0290050d",
   448 => x"0402f805",
   449 => x"0d8bb42d",
   450 => x"e008708b",
   451 => x"2a708106",
   452 => x"51525270",
   453 => x"802e9d38",
   454 => x"bbec0870",
   455 => x"8429bbf4",
   456 => x"057381ff",
   457 => x"06710c51",
   458 => x"51bbec08",
   459 => x"81118706",
   460 => x"bbec0c51",
   461 => x"800bbc94",
   462 => x"0c8ba72d",
   463 => x"8bae2d02",
   464 => x"88050d04",
   465 => x"02fc050d",
   466 => x"bbec518d",
   467 => x"aa2d8cd4",
   468 => x"2d8e8151",
   469 => x"8ba32d02",
   470 => x"84050d04",
   471 => x"bc9808bb",
   472 => x"c40c0402",
   473 => x"fc050d8e",
   474 => x"ed048bba",
   475 => x"2d80f651",
   476 => x"8cf12dbb",
   477 => x"c408f338",
   478 => x"80da518c",
   479 => x"f12dbbc4",
   480 => x"08e838bb",
   481 => x"c408ba84",
   482 => x"0cbbc408",
   483 => x"5184f02d",
   484 => x"0284050d",
   485 => x"0402ec05",
   486 => x"0d765480",
   487 => x"52870b88",
   488 => x"1580f52d",
   489 => x"56537472",
   490 => x"248338a0",
   491 => x"53725182",
   492 => x"f92d8112",
   493 => x"8b1580f5",
   494 => x"2d545272",
   495 => x"7225de38",
   496 => x"0294050d",
   497 => x"0402f005",
   498 => x"0dbc9808",
   499 => x"5481f82d",
   500 => x"800bbc9c",
   501 => x"0c730880",
   502 => x"2e818038",
   503 => x"820bbbd8",
   504 => x"0cbc9c08",
   505 => x"8f06bbd4",
   506 => x"0c730852",
   507 => x"71832e96",
   508 => x"38718326",
   509 => x"89387181",
   510 => x"2eaf3890",
   511 => x"c6047185",
   512 => x"2e9f3890",
   513 => x"c6048814",
   514 => x"80f52d84",
   515 => x"1508b5cc",
   516 => x"53545285",
   517 => x"fe2d7184",
   518 => x"29137008",
   519 => x"525290ca",
   520 => x"0473518f",
   521 => x"952d90c6",
   522 => x"04ba8008",
   523 => x"8815082c",
   524 => x"70810651",
   525 => x"5271802e",
   526 => x"8738b5d0",
   527 => x"5190c304",
   528 => x"b5d45185",
   529 => x"fe2d8414",
   530 => x"085185fe",
   531 => x"2dbc9c08",
   532 => x"8105bc9c",
   533 => x"0c8c1454",
   534 => x"8fd50402",
   535 => x"90050d04",
   536 => x"71bc980c",
   537 => x"8fc52dbc",
   538 => x"9c08ff05",
   539 => x"bca00c04",
   540 => x"02e8050d",
   541 => x"bc9808bc",
   542 => x"a4085755",
   543 => x"87518cf1",
   544 => x"2dbbc408",
   545 => x"812a7081",
   546 => x"06515271",
   547 => x"802ea038",
   548 => x"9196048b",
   549 => x"ba2d8751",
   550 => x"8cf12dbb",
   551 => x"c408f438",
   552 => x"ba840881",
   553 => x"3270ba84",
   554 => x"0c705252",
   555 => x"84f02d80",
   556 => x"fe518cf1",
   557 => x"2dbbc408",
   558 => x"802ea638",
   559 => x"ba840880",
   560 => x"2e913880",
   561 => x"0bba840c",
   562 => x"805184f0",
   563 => x"2d91d304",
   564 => x"8bba2d80",
   565 => x"fe518cf1",
   566 => x"2dbbc408",
   567 => x"f33886e2",
   568 => x"2dba8408",
   569 => x"903881fd",
   570 => x"518cf12d",
   571 => x"81fa518c",
   572 => x"f12d97a6",
   573 => x"0481f551",
   574 => x"8cf12dbb",
   575 => x"c408812a",
   576 => x"70810651",
   577 => x"5271802e",
   578 => x"af38bca0",
   579 => x"08527180",
   580 => x"2e8938ff",
   581 => x"12bca00c",
   582 => x"92b804bc",
   583 => x"9c0810bc",
   584 => x"9c080570",
   585 => x"84291651",
   586 => x"52881208",
   587 => x"802e8938",
   588 => x"ff518812",
   589 => x"0852712d",
   590 => x"81f2518c",
   591 => x"f12dbbc4",
   592 => x"08812a70",
   593 => x"81065152",
   594 => x"71802eb1",
   595 => x"38bc9c08",
   596 => x"ff11bca0",
   597 => x"08565353",
   598 => x"73722589",
   599 => x"388114bc",
   600 => x"a00c92fd",
   601 => x"04721013",
   602 => x"70842916",
   603 => x"51528812",
   604 => x"08802e89",
   605 => x"38fe5188",
   606 => x"12085271",
   607 => x"2d81fd51",
   608 => x"8cf12dbb",
   609 => x"c408812a",
   610 => x"70810651",
   611 => x"5271802e",
   612 => x"ad38bca0",
   613 => x"08802e89",
   614 => x"38800bbc",
   615 => x"a00c93be",
   616 => x"04bc9c08",
   617 => x"10bc9c08",
   618 => x"05708429",
   619 => x"16515288",
   620 => x"1208802e",
   621 => x"8938fd51",
   622 => x"88120852",
   623 => x"712d81fa",
   624 => x"518cf12d",
   625 => x"bbc40881",
   626 => x"2a708106",
   627 => x"51527180",
   628 => x"2eae38bc",
   629 => x"9c08ff11",
   630 => x"5452bca0",
   631 => x"08732588",
   632 => x"3872bca0",
   633 => x"0c948004",
   634 => x"71101270",
   635 => x"84291651",
   636 => x"52881208",
   637 => x"802e8938",
   638 => x"fc518812",
   639 => x"0852712d",
   640 => x"bca00870",
   641 => x"53547380",
   642 => x"2e8a388c",
   643 => x"15ff1555",
   644 => x"55948604",
   645 => x"820bbbd8",
   646 => x"0c718f06",
   647 => x"bbd40c81",
   648 => x"eb518cf1",
   649 => x"2dbbc408",
   650 => x"812a7081",
   651 => x"06515271",
   652 => x"802ead38",
   653 => x"7408852e",
   654 => x"098106a4",
   655 => x"38881580",
   656 => x"f52dff05",
   657 => x"52718816",
   658 => x"81b72d71",
   659 => x"982b5271",
   660 => x"80258838",
   661 => x"800b8816",
   662 => x"81b72d74",
   663 => x"518f952d",
   664 => x"81f4518c",
   665 => x"f12dbbc4",
   666 => x"08812a70",
   667 => x"81065152",
   668 => x"71802eb3",
   669 => x"38740885",
   670 => x"2e098106",
   671 => x"aa388815",
   672 => x"80f52d81",
   673 => x"05527188",
   674 => x"1681b72d",
   675 => x"7181ff06",
   676 => x"8b1680f5",
   677 => x"2d545272",
   678 => x"72278738",
   679 => x"72881681",
   680 => x"b72d7451",
   681 => x"8f952d80",
   682 => x"da518cf1",
   683 => x"2dbbc408",
   684 => x"812a7081",
   685 => x"06515271",
   686 => x"802e81a6",
   687 => x"38bc9808",
   688 => x"bca00855",
   689 => x"5373802e",
   690 => x"8a388c13",
   691 => x"ff155553",
   692 => x"95c50472",
   693 => x"08527182",
   694 => x"2ea63871",
   695 => x"82268938",
   696 => x"71812ea9",
   697 => x"3896e204",
   698 => x"71832eb1",
   699 => x"3871842e",
   700 => x"09810680",
   701 => x"ed388813",
   702 => x"085190e0",
   703 => x"2d96e204",
   704 => x"bca00851",
   705 => x"88130852",
   706 => x"712d96e2",
   707 => x"04810b88",
   708 => x"14082bba",
   709 => x"800832ba",
   710 => x"800c96b8",
   711 => x"04881380",
   712 => x"f52d8105",
   713 => x"8b1480f5",
   714 => x"2d535471",
   715 => x"74248338",
   716 => x"80547388",
   717 => x"1481b72d",
   718 => x"8fc52d96",
   719 => x"e2047508",
   720 => x"802ea238",
   721 => x"7508518c",
   722 => x"f12dbbc4",
   723 => x"08810652",
   724 => x"71802e8b",
   725 => x"38bca008",
   726 => x"51841608",
   727 => x"52712d88",
   728 => x"165675da",
   729 => x"38805480",
   730 => x"0bbbd80c",
   731 => x"738f06bb",
   732 => x"d40ca052",
   733 => x"73bca008",
   734 => x"2e098106",
   735 => x"9838bc9c",
   736 => x"08ff0574",
   737 => x"32700981",
   738 => x"05707207",
   739 => x"9f2a9171",
   740 => x"31515153",
   741 => x"53715182",
   742 => x"f92d8114",
   743 => x"548e7425",
   744 => x"c638ba84",
   745 => x"085271bb",
   746 => x"c40c0298",
   747 => x"050d0402",
   748 => x"f4050dd4",
   749 => x"5281ff72",
   750 => x"0c710853",
   751 => x"81ff720c",
   752 => x"72882b83",
   753 => x"fe800672",
   754 => x"087081ff",
   755 => x"06515253",
   756 => x"81ff720c",
   757 => x"72710788",
   758 => x"2b720870",
   759 => x"81ff0651",
   760 => x"525381ff",
   761 => x"720c7271",
   762 => x"07882b72",
   763 => x"087081ff",
   764 => x"067207bb",
   765 => x"c40c5253",
   766 => x"028c050d",
   767 => x"0402f405",
   768 => x"0d747671",
   769 => x"81ff06d4",
   770 => x"0c5353bc",
   771 => x"a8088538",
   772 => x"71892b52",
   773 => x"71982ad4",
   774 => x"0c71902a",
   775 => x"7081ff06",
   776 => x"d40c5171",
   777 => x"882a7081",
   778 => x"ff06d40c",
   779 => x"517181ff",
   780 => x"06d40c72",
   781 => x"902a7081",
   782 => x"ff06d40c",
   783 => x"51d40870",
   784 => x"81ff0651",
   785 => x"5182b8bf",
   786 => x"527081ff",
   787 => x"2e098106",
   788 => x"943881ff",
   789 => x"0bd40cd4",
   790 => x"087081ff",
   791 => x"06ff1454",
   792 => x"515171e5",
   793 => x"3870bbc4",
   794 => x"0c028c05",
   795 => x"0d0402fc",
   796 => x"050d81c7",
   797 => x"5181ff0b",
   798 => x"d40cff11",
   799 => x"51708025",
   800 => x"f4380284",
   801 => x"050d0402",
   802 => x"f4050d81",
   803 => x"ff0bd40c",
   804 => x"93538052",
   805 => x"87fc80c1",
   806 => x"5197fd2d",
   807 => x"bbc4088b",
   808 => x"3881ff0b",
   809 => x"d40c8153",
   810 => x"99b40498",
   811 => x"ee2dff13",
   812 => x"5372df38",
   813 => x"72bbc40c",
   814 => x"028c050d",
   815 => x"0402ec05",
   816 => x"0d810bbc",
   817 => x"a80c8454",
   818 => x"d008708f",
   819 => x"2a708106",
   820 => x"51515372",
   821 => x"f33872d0",
   822 => x"0c98ee2d",
   823 => x"b5d85185",
   824 => x"fe2dd008",
   825 => x"708f2a70",
   826 => x"81065151",
   827 => x"5372f338",
   828 => x"810bd00c",
   829 => x"b1538052",
   830 => x"84d480c0",
   831 => x"5197fd2d",
   832 => x"bbc40881",
   833 => x"2e933872",
   834 => x"822ebd38",
   835 => x"ff135372",
   836 => x"e538ff14",
   837 => x"5473ffb0",
   838 => x"3898ee2d",
   839 => x"83aa5284",
   840 => x"9c80c851",
   841 => x"97fd2dbb",
   842 => x"c408812e",
   843 => x"09810692",
   844 => x"3897af2d",
   845 => x"bbc40883",
   846 => x"ffff0653",
   847 => x"7283aa2e",
   848 => x"9d389987",
   849 => x"2d9ad904",
   850 => x"b5e45185",
   851 => x"fe2d8053",
   852 => x"9ca704b5",
   853 => x"fc5185fe",
   854 => x"2d80549b",
   855 => x"f90481ff",
   856 => x"0bd40cb1",
   857 => x"5498ee2d",
   858 => x"8fcf5380",
   859 => x"5287fc80",
   860 => x"f75197fd",
   861 => x"2dbbc408",
   862 => x"55bbc408",
   863 => x"812e0981",
   864 => x"069b3881",
   865 => x"ff0bd40c",
   866 => x"820a5284",
   867 => x"9c80e951",
   868 => x"97fd2dbb",
   869 => x"c408802e",
   870 => x"8d3898ee",
   871 => x"2dff1353",
   872 => x"72c9389b",
   873 => x"ec0481ff",
   874 => x"0bd40cbb",
   875 => x"c4085287",
   876 => x"fc80fa51",
   877 => x"97fd2dbb",
   878 => x"c408b138",
   879 => x"81ff0bd4",
   880 => x"0cd40853",
   881 => x"81ff0bd4",
   882 => x"0c81ff0b",
   883 => x"d40c81ff",
   884 => x"0bd40c81",
   885 => x"ff0bd40c",
   886 => x"72862a70",
   887 => x"81067656",
   888 => x"51537295",
   889 => x"38bbc408",
   890 => x"549bf904",
   891 => x"73822efe",
   892 => x"e238ff14",
   893 => x"5473feed",
   894 => x"3873bca8",
   895 => x"0c738b38",
   896 => x"815287fc",
   897 => x"80d05197",
   898 => x"fd2d81ff",
   899 => x"0bd40cd0",
   900 => x"08708f2a",
   901 => x"70810651",
   902 => x"515372f3",
   903 => x"3872d00c",
   904 => x"81ff0bd4",
   905 => x"0c815372",
   906 => x"bbc40c02",
   907 => x"94050d04",
   908 => x"02e8050d",
   909 => x"78558056",
   910 => x"81ff0bd4",
   911 => x"0cd00870",
   912 => x"8f2a7081",
   913 => x"06515153",
   914 => x"72f33882",
   915 => x"810bd00c",
   916 => x"81ff0bd4",
   917 => x"0c775287",
   918 => x"fc80d151",
   919 => x"97fd2d80",
   920 => x"dbc6df54",
   921 => x"bbc40880",
   922 => x"2e8a38b6",
   923 => x"9c5185fe",
   924 => x"2d9dc704",
   925 => x"81ff0bd4",
   926 => x"0cd40870",
   927 => x"81ff0651",
   928 => x"537281fe",
   929 => x"2e098106",
   930 => x"9d3880ff",
   931 => x"5397af2d",
   932 => x"bbc40875",
   933 => x"70840557",
   934 => x"0cff1353",
   935 => x"728025ed",
   936 => x"3881569d",
   937 => x"ac04ff14",
   938 => x"5473c938",
   939 => x"81ff0bd4",
   940 => x"0c81ff0b",
   941 => x"d40cd008",
   942 => x"708f2a70",
   943 => x"81065151",
   944 => x"5372f338",
   945 => x"72d00c75",
   946 => x"bbc40c02",
   947 => x"98050d04",
   948 => x"02e8050d",
   949 => x"77797b58",
   950 => x"55558053",
   951 => x"727625a3",
   952 => x"38747081",
   953 => x"055680f5",
   954 => x"2d747081",
   955 => x"055680f5",
   956 => x"2d525271",
   957 => x"712e8638",
   958 => x"81519e85",
   959 => x"04811353",
   960 => x"9ddc0480",
   961 => x"5170bbc4",
   962 => x"0c029805",
   963 => x"0d0402ec",
   964 => x"050d7655",
   965 => x"74802ebe",
   966 => x"389a1580",
   967 => x"e02d51ab",
   968 => x"ce2dbbc4",
   969 => x"08bbc408",
   970 => x"80c2dc0c",
   971 => x"bbc40854",
   972 => x"5480c2b8",
   973 => x"08802e99",
   974 => x"38941580",
   975 => x"e02d51ab",
   976 => x"ce2dbbc4",
   977 => x"08902b83",
   978 => x"fff00a06",
   979 => x"70750751",
   980 => x"537280c2",
   981 => x"dc0c80c2",
   982 => x"dc085372",
   983 => x"802e9d38",
   984 => x"80c2b008",
   985 => x"fe147129",
   986 => x"80c2c408",
   987 => x"0580c2e0",
   988 => x"0c70842b",
   989 => x"80c2bc0c",
   990 => x"549faa04",
   991 => x"80c2c808",
   992 => x"80c2dc0c",
   993 => x"80c2cc08",
   994 => x"80c2e00c",
   995 => x"80c2b808",
   996 => x"802e8b38",
   997 => x"80c2b008",
   998 => x"842b539f",
   999 => x"a50480c2",
  1000 => x"d008842b",
  1001 => x"537280c2",
  1002 => x"bc0c0294",
  1003 => x"050d0402",
  1004 => x"d8050d80",
  1005 => x"0b80c2b8",
  1006 => x"0c845499",
  1007 => x"bd2dbbc4",
  1008 => x"08802e95",
  1009 => x"38bcac52",
  1010 => x"80519cb0",
  1011 => x"2dbbc408",
  1012 => x"802e8638",
  1013 => x"fe549fe1",
  1014 => x"04ff1454",
  1015 => x"738024db",
  1016 => x"38738c38",
  1017 => x"b6ac5185",
  1018 => x"fe2d7355",
  1019 => x"a5870480",
  1020 => x"56810b80",
  1021 => x"c2e40c88",
  1022 => x"53b6c052",
  1023 => x"bce2519d",
  1024 => x"d02dbbc4",
  1025 => x"08762e09",
  1026 => x"81068838",
  1027 => x"bbc40880",
  1028 => x"c2e40c88",
  1029 => x"53b6cc52",
  1030 => x"bcfe519d",
  1031 => x"d02dbbc4",
  1032 => x"088838bb",
  1033 => x"c40880c2",
  1034 => x"e40c80c2",
  1035 => x"e408802e",
  1036 => x"80f838bf",
  1037 => x"f20b80f5",
  1038 => x"2dbff30b",
  1039 => x"80f52d71",
  1040 => x"982b7190",
  1041 => x"2b07bff4",
  1042 => x"0b80f52d",
  1043 => x"70882b72",
  1044 => x"07bff50b",
  1045 => x"80f52d71",
  1046 => x"0780c0aa",
  1047 => x"0b80f52d",
  1048 => x"80c0ab0b",
  1049 => x"80f52d71",
  1050 => x"882b0753",
  1051 => x"5f54525a",
  1052 => x"56575573",
  1053 => x"81abaa2e",
  1054 => x"0981068d",
  1055 => x"387551ab",
  1056 => x"9e2dbbc4",
  1057 => x"0856a196",
  1058 => x"047382d4",
  1059 => x"d52e8738",
  1060 => x"b6d851a1",
  1061 => x"d804bcac",
  1062 => x"5275519c",
  1063 => x"b02dbbc4",
  1064 => x"0855bbc4",
  1065 => x"08802e83",
  1066 => x"de388853",
  1067 => x"b6cc52bc",
  1068 => x"fe519dd0",
  1069 => x"2dbbc408",
  1070 => x"8a38810b",
  1071 => x"80c2b80c",
  1072 => x"a1de0488",
  1073 => x"53b6c052",
  1074 => x"bce2519d",
  1075 => x"d02dbbc4",
  1076 => x"08802e8a",
  1077 => x"38b6ec51",
  1078 => x"85fe2da2",
  1079 => x"ba0480c0",
  1080 => x"aa0b80f5",
  1081 => x"2d547380",
  1082 => x"d52e0981",
  1083 => x"0680cb38",
  1084 => x"80c0ab0b",
  1085 => x"80f52d54",
  1086 => x"7381aa2e",
  1087 => x"098106ba",
  1088 => x"38800bbc",
  1089 => x"ac0b80f5",
  1090 => x"2d565474",
  1091 => x"81e92e83",
  1092 => x"38815474",
  1093 => x"81eb2e8c",
  1094 => x"38805573",
  1095 => x"752e0981",
  1096 => x"0682e438",
  1097 => x"bcb70b80",
  1098 => x"f52d5574",
  1099 => x"8d38bcb8",
  1100 => x"0b80f52d",
  1101 => x"5473822e",
  1102 => x"86388055",
  1103 => x"a58704bc",
  1104 => x"b90b80f5",
  1105 => x"2d7080c2",
  1106 => x"b00cff05",
  1107 => x"80c2b40c",
  1108 => x"bcba0b80",
  1109 => x"f52dbcbb",
  1110 => x"0b80f52d",
  1111 => x"58760577",
  1112 => x"82802905",
  1113 => x"7080c2c0",
  1114 => x"0cbcbc0b",
  1115 => x"80f52d70",
  1116 => x"80c2d40c",
  1117 => x"80c2b808",
  1118 => x"59575876",
  1119 => x"802e81ac",
  1120 => x"388853b6",
  1121 => x"cc52bcfe",
  1122 => x"519dd02d",
  1123 => x"bbc40881",
  1124 => x"f63880c2",
  1125 => x"b0087084",
  1126 => x"2b80c2bc",
  1127 => x"0c7080c2",
  1128 => x"d00cbcd1",
  1129 => x"0b80f52d",
  1130 => x"bcd00b80",
  1131 => x"f52d7182",
  1132 => x"802905bc",
  1133 => x"d20b80f5",
  1134 => x"2d708480",
  1135 => x"802912bc",
  1136 => x"d30b80f5",
  1137 => x"2d708180",
  1138 => x"0a291270",
  1139 => x"80c2d80c",
  1140 => x"80c2d408",
  1141 => x"712980c2",
  1142 => x"c0080570",
  1143 => x"80c2c40c",
  1144 => x"bcd90b80",
  1145 => x"f52dbcd8",
  1146 => x"0b80f52d",
  1147 => x"71828029",
  1148 => x"05bcda0b",
  1149 => x"80f52d70",
  1150 => x"84808029",
  1151 => x"12bcdb0b",
  1152 => x"80f52d70",
  1153 => x"982b81f0",
  1154 => x"0a067205",
  1155 => x"7080c2c8",
  1156 => x"0cfe117e",
  1157 => x"29770580",
  1158 => x"c2cc0c52",
  1159 => x"59524354",
  1160 => x"5e515259",
  1161 => x"525d5759",
  1162 => x"57a58004",
  1163 => x"bcbe0b80",
  1164 => x"f52dbcbd",
  1165 => x"0b80f52d",
  1166 => x"71828029",
  1167 => x"057080c2",
  1168 => x"bc0c70a0",
  1169 => x"2983ff05",
  1170 => x"70892a70",
  1171 => x"80c2d00c",
  1172 => x"bcc30b80",
  1173 => x"f52dbcc2",
  1174 => x"0b80f52d",
  1175 => x"71828029",
  1176 => x"057080c2",
  1177 => x"d80c7b71",
  1178 => x"291e7080",
  1179 => x"c2cc0c7d",
  1180 => x"80c2c80c",
  1181 => x"730580c2",
  1182 => x"c40c555e",
  1183 => x"51515555",
  1184 => x"80519e8e",
  1185 => x"2d815574",
  1186 => x"bbc40c02",
  1187 => x"a8050d04",
  1188 => x"02ec050d",
  1189 => x"7670872c",
  1190 => x"7180ff06",
  1191 => x"55565480",
  1192 => x"c2b8088a",
  1193 => x"3873882c",
  1194 => x"7481ff06",
  1195 => x"5455bcac",
  1196 => x"5280c2c0",
  1197 => x"0815519c",
  1198 => x"b02dbbc4",
  1199 => x"0854bbc4",
  1200 => x"08802eb4",
  1201 => x"3880c2b8",
  1202 => x"08802e98",
  1203 => x"38728429",
  1204 => x"bcac0570",
  1205 => x"085253ab",
  1206 => x"9e2dbbc4",
  1207 => x"08f00a06",
  1208 => x"53a5f604",
  1209 => x"7210bcac",
  1210 => x"057080e0",
  1211 => x"2d5253ab",
  1212 => x"ce2dbbc4",
  1213 => x"08537254",
  1214 => x"73bbc40c",
  1215 => x"0294050d",
  1216 => x"0402e005",
  1217 => x"0d797084",
  1218 => x"2c80c2e0",
  1219 => x"0805718f",
  1220 => x"06525553",
  1221 => x"728938bc",
  1222 => x"ac527351",
  1223 => x"9cb02d72",
  1224 => x"a029bcac",
  1225 => x"05548074",
  1226 => x"80f52d56",
  1227 => x"5374732e",
  1228 => x"83388153",
  1229 => x"7481e52e",
  1230 => x"81f13881",
  1231 => x"70740654",
  1232 => x"5872802e",
  1233 => x"81e5388b",
  1234 => x"1480f52d",
  1235 => x"70832a79",
  1236 => x"06585676",
  1237 => x"9938ba88",
  1238 => x"08537289",
  1239 => x"387280c0",
  1240 => x"ac0b81b7",
  1241 => x"2d76ba88",
  1242 => x"0c7353a8",
  1243 => x"ad04758f",
  1244 => x"2e098106",
  1245 => x"81b53874",
  1246 => x"9f068d29",
  1247 => x"80c09f11",
  1248 => x"51538114",
  1249 => x"80f52d73",
  1250 => x"70810555",
  1251 => x"81b72d83",
  1252 => x"1480f52d",
  1253 => x"73708105",
  1254 => x"5581b72d",
  1255 => x"851480f5",
  1256 => x"2d737081",
  1257 => x"055581b7",
  1258 => x"2d871480",
  1259 => x"f52d7370",
  1260 => x"81055581",
  1261 => x"b72d8914",
  1262 => x"80f52d73",
  1263 => x"70810555",
  1264 => x"81b72d8e",
  1265 => x"1480f52d",
  1266 => x"73708105",
  1267 => x"5581b72d",
  1268 => x"901480f5",
  1269 => x"2d737081",
  1270 => x"055581b7",
  1271 => x"2d921480",
  1272 => x"f52d7370",
  1273 => x"81055581",
  1274 => x"b72d9414",
  1275 => x"80f52d73",
  1276 => x"70810555",
  1277 => x"81b72d96",
  1278 => x"1480f52d",
  1279 => x"73708105",
  1280 => x"5581b72d",
  1281 => x"981480f5",
  1282 => x"2d737081",
  1283 => x"055581b7",
  1284 => x"2d9c1480",
  1285 => x"f52d7370",
  1286 => x"81055581",
  1287 => x"b72d9e14",
  1288 => x"80f52d73",
  1289 => x"81b72d77",
  1290 => x"ba880c80",
  1291 => x"5372bbc4",
  1292 => x"0c02a005",
  1293 => x"0d0402cc",
  1294 => x"050d7e60",
  1295 => x"5e5a800b",
  1296 => x"80c2dc08",
  1297 => x"80c2e008",
  1298 => x"595c5680",
  1299 => x"5880c2bc",
  1300 => x"08782e81",
  1301 => x"b038778f",
  1302 => x"06a01757",
  1303 => x"54738f38",
  1304 => x"bcac5276",
  1305 => x"51811757",
  1306 => x"9cb02dbc",
  1307 => x"ac568076",
  1308 => x"80f52d56",
  1309 => x"5474742e",
  1310 => x"83388154",
  1311 => x"7481e52e",
  1312 => x"80f73881",
  1313 => x"70750655",
  1314 => x"5c73802e",
  1315 => x"80eb388b",
  1316 => x"1680f52d",
  1317 => x"98065978",
  1318 => x"80df388b",
  1319 => x"537c5275",
  1320 => x"519dd02d",
  1321 => x"bbc40880",
  1322 => x"d0389c16",
  1323 => x"0851ab9e",
  1324 => x"2dbbc408",
  1325 => x"841b0c9a",
  1326 => x"1680e02d",
  1327 => x"51abce2d",
  1328 => x"bbc408bb",
  1329 => x"c408881c",
  1330 => x"0cbbc408",
  1331 => x"555580c2",
  1332 => x"b808802e",
  1333 => x"98389416",
  1334 => x"80e02d51",
  1335 => x"abce2dbb",
  1336 => x"c408902b",
  1337 => x"83fff00a",
  1338 => x"06701651",
  1339 => x"5473881b",
  1340 => x"0c787a0c",
  1341 => x"7b54aabe",
  1342 => x"04811858",
  1343 => x"80c2bc08",
  1344 => x"7826fed2",
  1345 => x"3880c2b8",
  1346 => x"08802eb0",
  1347 => x"387a51a5",
  1348 => x"902dbbc4",
  1349 => x"08bbc408",
  1350 => x"80ffffff",
  1351 => x"f806555b",
  1352 => x"7380ffff",
  1353 => x"fff82e94",
  1354 => x"38bbc408",
  1355 => x"fe0580c2",
  1356 => x"b0082980",
  1357 => x"c2c40805",
  1358 => x"57a8cb04",
  1359 => x"805473bb",
  1360 => x"c40c02b4",
  1361 => x"050d0402",
  1362 => x"f4050d74",
  1363 => x"70088105",
  1364 => x"710c7008",
  1365 => x"80c2b408",
  1366 => x"06535371",
  1367 => x"8e388813",
  1368 => x"0851a590",
  1369 => x"2dbbc408",
  1370 => x"88140c81",
  1371 => x"0bbbc40c",
  1372 => x"028c050d",
  1373 => x"0402f005",
  1374 => x"0d758811",
  1375 => x"08fe0580",
  1376 => x"c2b00829",
  1377 => x"80c2c408",
  1378 => x"11720880",
  1379 => x"c2b40806",
  1380 => x"05795553",
  1381 => x"54549cb0",
  1382 => x"2d029005",
  1383 => x"0d0402f4",
  1384 => x"050d7470",
  1385 => x"882a83fe",
  1386 => x"80067072",
  1387 => x"982a0772",
  1388 => x"882b87fc",
  1389 => x"80800673",
  1390 => x"982b81f0",
  1391 => x"0a067173",
  1392 => x"0707bbc4",
  1393 => x"0c565153",
  1394 => x"51028c05",
  1395 => x"0d0402f8",
  1396 => x"050d028e",
  1397 => x"0580f52d",
  1398 => x"74882b07",
  1399 => x"7083ffff",
  1400 => x"06bbc40c",
  1401 => x"51028805",
  1402 => x"0d0402f4",
  1403 => x"050d7476",
  1404 => x"78535452",
  1405 => x"80712597",
  1406 => x"38727081",
  1407 => x"055480f5",
  1408 => x"2d727081",
  1409 => x"055481b7",
  1410 => x"2dff1151",
  1411 => x"70eb3880",
  1412 => x"7281b72d",
  1413 => x"028c050d",
  1414 => x"0402e805",
  1415 => x"0d775680",
  1416 => x"70565473",
  1417 => x"7624b338",
  1418 => x"80c2bc08",
  1419 => x"742eab38",
  1420 => x"7351a681",
  1421 => x"2dbbc408",
  1422 => x"bbc40809",
  1423 => x"810570bb",
  1424 => x"c408079f",
  1425 => x"2a770581",
  1426 => x"17575753",
  1427 => x"53747624",
  1428 => x"893880c2",
  1429 => x"bc087426",
  1430 => x"d73872bb",
  1431 => x"c40c0298",
  1432 => x"050d0402",
  1433 => x"f0050dbb",
  1434 => x"c0081651",
  1435 => x"ac992dbb",
  1436 => x"c408802e",
  1437 => x"9e388b53",
  1438 => x"bbc40852",
  1439 => x"80c0ac51",
  1440 => x"abea2d80",
  1441 => x"c2e80854",
  1442 => x"73802e87",
  1443 => x"3880c0ac",
  1444 => x"51732d02",
  1445 => x"90050d04",
  1446 => x"02dc050d",
  1447 => x"80705a55",
  1448 => x"74bbc008",
  1449 => x"25b13880",
  1450 => x"c2bc0875",
  1451 => x"2ea93878",
  1452 => x"51a6812d",
  1453 => x"bbc40809",
  1454 => x"810570bb",
  1455 => x"c408079f",
  1456 => x"2a760581",
  1457 => x"1b5b5654",
  1458 => x"74bbc008",
  1459 => x"25893880",
  1460 => x"c2bc0879",
  1461 => x"26d93880",
  1462 => x"557880c2",
  1463 => x"bc082781",
  1464 => x"d4387851",
  1465 => x"a6812dbb",
  1466 => x"c408802e",
  1467 => x"81a838bb",
  1468 => x"c4088b05",
  1469 => x"80f52d70",
  1470 => x"842a7081",
  1471 => x"06771078",
  1472 => x"842b80c0",
  1473 => x"ac0b80f5",
  1474 => x"2d5c5c53",
  1475 => x"51555673",
  1476 => x"802e80c9",
  1477 => x"38741682",
  1478 => x"2bafd90b",
  1479 => x"ba94120c",
  1480 => x"54777531",
  1481 => x"1080c2ec",
  1482 => x"11555690",
  1483 => x"74708105",
  1484 => x"5681b72d",
  1485 => x"a07481b7",
  1486 => x"2d7681ff",
  1487 => x"06811658",
  1488 => x"5473802e",
  1489 => x"8a389c53",
  1490 => x"80c0ac52",
  1491 => x"aed5048b",
  1492 => x"53bbc408",
  1493 => x"5280c2ee",
  1494 => x"1651af8e",
  1495 => x"04741682",
  1496 => x"2bace30b",
  1497 => x"ba94120c",
  1498 => x"547681ff",
  1499 => x"06811658",
  1500 => x"5473802e",
  1501 => x"8a389c53",
  1502 => x"80c0ac52",
  1503 => x"af85048b",
  1504 => x"53bbc408",
  1505 => x"52777531",
  1506 => x"1080c2ec",
  1507 => x"05517655",
  1508 => x"abea2daf",
  1509 => x"aa047490",
  1510 => x"29753170",
  1511 => x"1080c2ec",
  1512 => x"055154bb",
  1513 => x"c4087481",
  1514 => x"b72d8119",
  1515 => x"59748b24",
  1516 => x"a338add9",
  1517 => x"04749029",
  1518 => x"75317010",
  1519 => x"80c2ec05",
  1520 => x"8c773157",
  1521 => x"51548074",
  1522 => x"81b72d9e",
  1523 => x"14ff1656",
  1524 => x"5474f338",
  1525 => x"02a4050d",
  1526 => x"0402fc05",
  1527 => x"0dbbc008",
  1528 => x"1351ac99",
  1529 => x"2dbbc408",
  1530 => x"802e8838",
  1531 => x"bbc40851",
  1532 => x"9e8e2d80",
  1533 => x"0bbbc00c",
  1534 => x"ad982d8f",
  1535 => x"c52d0284",
  1536 => x"050d0402",
  1537 => x"fc050d72",
  1538 => x"5170fd2e",
  1539 => x"ad3870fd",
  1540 => x"248a3870",
  1541 => x"fc2e80c4",
  1542 => x"38b0e404",
  1543 => x"70fe2eb1",
  1544 => x"3870ff2e",
  1545 => x"098106bc",
  1546 => x"38bbc008",
  1547 => x"5170802e",
  1548 => x"b338ff11",
  1549 => x"bbc00cb0",
  1550 => x"e404bbc0",
  1551 => x"08f00570",
  1552 => x"bbc00c51",
  1553 => x"7080259c",
  1554 => x"38800bbb",
  1555 => x"c00cb0e4",
  1556 => x"04bbc008",
  1557 => x"8105bbc0",
  1558 => x"0cb0e404",
  1559 => x"bbc00890",
  1560 => x"05bbc00c",
  1561 => x"ad982d8f",
  1562 => x"c52d0284",
  1563 => x"050d0402",
  1564 => x"fc050d80",
  1565 => x"0bbbc00c",
  1566 => x"ad982d8e",
  1567 => x"dc2dbbc4",
  1568 => x"08bbb00c",
  1569 => x"ba8c5190",
  1570 => x"e02d0284",
  1571 => x"050d0471",
  1572 => x"80c2e80c",
  1573 => x"04000000",
  1574 => x"00ffffff",
  1575 => x"ff00ffff",
  1576 => x"ffff00ff",
  1577 => x"ffffff00",
  1578 => x"52657365",
  1579 => x"74000000",
  1580 => x"43617267",
  1581 => x"61722044",
  1582 => x"6973636f",
  1583 => x"2f43696e",
  1584 => x"74612010",
  1585 => x"00000000",
  1586 => x"45786974",
  1587 => x"00000000",
  1588 => x"43617267",
  1589 => x"61206465",
  1590 => x"2043696e",
  1591 => x"74612052",
  1592 => x"61706964",
  1593 => x"61000000",
  1594 => x"43617267",
  1595 => x"61206465",
  1596 => x"2043696e",
  1597 => x"7461204e",
  1598 => x"6f726d61",
  1599 => x"6c000000",
  1600 => x"53706563",
  1601 => x"7472756d",
  1602 => x"20313238",
  1603 => x"4b000000",
  1604 => x"50656e74",
  1605 => x"61676f6e",
  1606 => x"20313032",
  1607 => x"344b0000",
  1608 => x"50726f66",
  1609 => x"69203130",
  1610 => x"32344b00",
  1611 => x"53706563",
  1612 => x"7472756d",
  1613 => x"2034384b",
  1614 => x"00000000",
  1615 => x"53706563",
  1616 => x"7472756d",
  1617 => x"202b3241",
  1618 => x"2f2b3300",
  1619 => x"554c412d",
  1620 => x"34380000",
  1621 => x"554c412d",
  1622 => x"31323800",
  1623 => x"50656e74",
  1624 => x"61676f6e",
  1625 => x"00000000",
  1626 => x"556c612b",
  1627 => x"20262054",
  1628 => x"696d6578",
  1629 => x"00000000",
  1630 => x"4e6f726d",
  1631 => x"616c0000",
  1632 => x"47656e65",
  1633 => x"72616c20",
  1634 => x"536f756e",
  1635 => x"6420324d",
  1636 => x"42000000",
  1637 => x"47656e65",
  1638 => x"72616c20",
  1639 => x"536f756e",
  1640 => x"64204465",
  1641 => x"73616374",
  1642 => x"69766164",
  1643 => x"6f000000",
  1644 => x"4d4d4320",
  1645 => x"43617264",
  1646 => x"206f6666",
  1647 => x"00000000",
  1648 => x"6469764d",
  1649 => x"4d430000",
  1650 => x"5a584d4d",
  1651 => x"43000000",
  1652 => x"4a6f7920",
  1653 => x"323a2053",
  1654 => x"696e636c",
  1655 => x"61697220",
  1656 => x"49000000",
  1657 => x"4a6f7920",
  1658 => x"323a2053",
  1659 => x"696e636c",
  1660 => x"61697220",
  1661 => x"49490000",
  1662 => x"4a6f7920",
  1663 => x"323a204b",
  1664 => x"656d7374",
  1665 => x"6f6e0000",
  1666 => x"4a6f7920",
  1667 => x"323a2043",
  1668 => x"7572736f",
  1669 => x"72000000",
  1670 => x"4a6f7920",
  1671 => x"313a2053",
  1672 => x"696e636c",
  1673 => x"61697220",
  1674 => x"49000000",
  1675 => x"4a6f7920",
  1676 => x"313a2053",
  1677 => x"696e636c",
  1678 => x"61697220",
  1679 => x"49490000",
  1680 => x"4a6f7920",
  1681 => x"313a204b",
  1682 => x"656d7374",
  1683 => x"6f6e0000",
  1684 => x"4a6f7920",
  1685 => x"313a2043",
  1686 => x"7572736f",
  1687 => x"72000000",
  1688 => x"5363616e",
  1689 => x"6c696e65",
  1690 => x"73204e6f",
  1691 => x"6e650000",
  1692 => x"5363616e",
  1693 => x"6c696e65",
  1694 => x"73204352",
  1695 => x"54203235",
  1696 => x"25000000",
  1697 => x"5363616e",
  1698 => x"6c696e65",
  1699 => x"73204352",
  1700 => x"54203530",
  1701 => x"25000000",
  1702 => x"5363616e",
  1703 => x"6c696e65",
  1704 => x"73204352",
  1705 => x"54203735",
  1706 => x"25000000",
  1707 => x"43617267",
  1708 => x"61204661",
  1709 => x"6c6c6964",
  1710 => x"61000000",
  1711 => x"4f4b0000",
  1712 => x"53504543",
  1713 => x"5452554d",
  1714 => x"44415400",
  1715 => x"16200000",
  1716 => x"14200000",
  1717 => x"15200000",
  1718 => x"53442069",
  1719 => x"6e69742e",
  1720 => x"2e2e0a00",
  1721 => x"53442063",
  1722 => x"61726420",
  1723 => x"72657365",
  1724 => x"74206661",
  1725 => x"696c6564",
  1726 => x"210a0000",
  1727 => x"53444843",
  1728 => x"20657272",
  1729 => x"6f72210a",
  1730 => x"00000000",
  1731 => x"57726974",
  1732 => x"65206661",
  1733 => x"696c6564",
  1734 => x"0a000000",
  1735 => x"52656164",
  1736 => x"20666169",
  1737 => x"6c65640a",
  1738 => x"00000000",
  1739 => x"43617264",
  1740 => x"20696e69",
  1741 => x"74206661",
  1742 => x"696c6564",
  1743 => x"0a000000",
  1744 => x"46415431",
  1745 => x"36202020",
  1746 => x"00000000",
  1747 => x"46415433",
  1748 => x"32202020",
  1749 => x"00000000",
  1750 => x"4e6f2070",
  1751 => x"61727469",
  1752 => x"74696f6e",
  1753 => x"20736967",
  1754 => x"0a000000",
  1755 => x"42616420",
  1756 => x"70617274",
  1757 => x"0a000000",
  1758 => x"4261636b",
  1759 => x"00000000",
  1760 => x"00000002",
  1761 => x"00000002",
  1762 => x"000018a8",
  1763 => x"0000034e",
  1764 => x"00000003",
  1765 => x"00001c84",
  1766 => x"00000004",
  1767 => x"00000003",
  1768 => x"00001c74",
  1769 => x"00000005",
  1770 => x"00000003",
  1771 => x"00001c64",
  1772 => x"00000005",
  1773 => x"00000003",
  1774 => x"00001c58",
  1775 => x"00000003",
  1776 => x"00000003",
  1777 => x"00001c50",
  1778 => x"00000002",
  1779 => x"00000003",
  1780 => x"00001c48",
  1781 => x"00000002",
  1782 => x"00000003",
  1783 => x"00001c3c",
  1784 => x"00000003",
  1785 => x"00000003",
  1786 => x"00001c28",
  1787 => x"00000005",
  1788 => x"00000003",
  1789 => x"00001c20",
  1790 => x"00000002",
  1791 => x"00000002",
  1792 => x"000018b0",
  1793 => x"0000186f",
  1794 => x"00000002",
  1795 => x"000018c8",
  1796 => x"00000763",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"00000000",
  1800 => x"000018d0",
  1801 => x"000018e8",
  1802 => x"00001900",
  1803 => x"00001910",
  1804 => x"00001920",
  1805 => x"0000192c",
  1806 => x"0000193c",
  1807 => x"0000194c",
  1808 => x"00001954",
  1809 => x"0000195c",
  1810 => x"00001968",
  1811 => x"00001978",
  1812 => x"00001980",
  1813 => x"00001994",
  1814 => x"000019b0",
  1815 => x"000019c0",
  1816 => x"000019c8",
  1817 => x"000019d0",
  1818 => x"000019e4",
  1819 => x"000019f8",
  1820 => x"00001a08",
  1821 => x"00001a18",
  1822 => x"00001a2c",
  1823 => x"00001a40",
  1824 => x"00001a50",
  1825 => x"00001a60",
  1826 => x"00001a70",
  1827 => x"00001a84",
  1828 => x"00001a98",
  1829 => x"00000004",
  1830 => x"00001aac",
  1831 => x"00001c94",
  1832 => x"00000004",
  1833 => x"00001abc",
  1834 => x"00001b84",
  1835 => x"00000000",
  1836 => x"00000000",
  1837 => x"00000000",
  1838 => x"00000000",
  1839 => x"00000000",
  1840 => x"00000000",
  1841 => x"00000000",
  1842 => x"00000000",
  1843 => x"00000000",
  1844 => x"00000000",
  1845 => x"00000000",
  1846 => x"00000000",
  1847 => x"00000000",
  1848 => x"00000000",
  1849 => x"00000000",
  1850 => x"00000000",
  1851 => x"00000000",
  1852 => x"00000000",
  1853 => x"00000000",
  1854 => x"00000000",
  1855 => x"00000000",
  1856 => x"00000000",
  1857 => x"00000000",
  1858 => x"00000000",
  1859 => x"00000002",
  1860 => x"0000216c",
  1861 => x"00001663",
  1862 => x"00000002",
  1863 => x"0000218a",
  1864 => x"00001663",
  1865 => x"00000002",
  1866 => x"000021a8",
  1867 => x"00001663",
  1868 => x"00000002",
  1869 => x"000021c6",
  1870 => x"00001663",
  1871 => x"00000002",
  1872 => x"000021e4",
  1873 => x"00001663",
  1874 => x"00000002",
  1875 => x"00002202",
  1876 => x"00001663",
  1877 => x"00000002",
  1878 => x"00002220",
  1879 => x"00001663",
  1880 => x"00000002",
  1881 => x"0000223e",
  1882 => x"00001663",
  1883 => x"00000002",
  1884 => x"0000225c",
  1885 => x"00001663",
  1886 => x"00000002",
  1887 => x"0000227a",
  1888 => x"00001663",
  1889 => x"00000002",
  1890 => x"00002298",
  1891 => x"00001663",
  1892 => x"00000002",
  1893 => x"000022b6",
  1894 => x"00001663",
  1895 => x"00000002",
  1896 => x"000022d4",
  1897 => x"00001663",
  1898 => x"00000004",
  1899 => x"00001b78",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"00001803",
  1904 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

